
.param mc_mm_switch=0
.param mc_pr_switch=0
.include /media/ASIC/caravel_FlexRV32/dependencies/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /media/ASIC/caravel_FlexRV32/dependencies/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /media/ASIC/caravel_FlexRV32/dependencies/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /media/ASIC/caravel_FlexRV32/dependencies/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice
.include /media/ASIC/caravel_FlexRV32/dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
