* NGSPICE file created from rv_alu1.ext - technology: sky130A


X_432_ _109_ VSS VSS VCC VCC o_op1[9] sky130_fd_sc_hd__buf_2
X_501_ i_reg2_data[11] imm_i\[11\] _142_ VSS VSS VCC VCC _145_ sky130_fd_sc_hd__mux2_1
X_981_ clknet_3_7__leaf_i_clk _040_ VSS VSS VCC VCC o_to_trap sky130_fd_sc_hd__dfxtp_2
X_415_ _100_ VSS VSS VCC VCC o_op1[1] sky130_fd_sc_hd__buf_2
X_964_ clknet_3_5__leaf_i_clk _023_ VSS VSS VCC VCC o_funct3[1] sky130_fd_sc_hd__dfxtp_2
X_895_ _407_ VSS VSS VCC VCC _053_ sky130_fd_sc_hd__clkbuf_1
X_680_ i_rs1[2] o_rs1[2] _282_ VSS VSS VCC VCC _285_ sky130_fd_sc_hd__mux2_1
X_878_ i_pc_next[5] o_pc_next[5] _390_ VSS VSS VCC VCC _399_ sky130_fd_sc_hd__mux2_1
X_947_ clknet_3_0__leaf_i_clk _006_ VSS VSS VCC VCC op1_sel sky130_fd_sc_hd__dfxtp_2
X_801_ _288_ VSS VSS VCC VCC _354_ sky130_fd_sc_hd__clkbuf_2
X_732_ _315_ VSS VSS VCC VCC _079_ sky130_fd_sc_hd__clkbuf_1
X_663_ imm_i\[15\] _271_ VSS VSS VCC VCC _272_ sky130_fd_sc_hd__or2_1
X_594_ _174_ _208_ _210_ VSS VSS VCC VCC _211_ sky130_fd_sc_hd__a21oi_1
X_715_ i_imm_i[0] imm_i\[0\] _306_ VSS VSS VCC VCC _307_ sky130_fd_sc_hd__mux2_1
X_646_ o_pc[13] i_reg1_data[13] _168_ VSS VSS VCC VCC _257_ sky130_fd_sc_hd__mux2_1
X_577_ o_pc[5] i_reg1_data[5] inst_jalr VSS VSS VCC VCC _196_ sky130_fd_sc_hd__mux2_1
X_500_ _144_ VSS VSS VCC VCC o_op2[10] sky130_fd_sc_hd__buf_2
X_431_ i_reg1_data[9] o_pc[9] _102_ VSS VSS VCC VCC _109_ sky130_fd_sc_hd__mux2_1
X_629_ _225_ imm_i\[11\] _241_ VSS VSS VCC VCC _242_ sky130_fd_sc_hd__and3_1
X_980_ clknet_3_3__leaf_i_clk _039_ VSS VSS VCC VCC o_pc[15] sky130_fd_sc_hd__dfxtp_2
X_414_ i_reg1_data[1] o_pc[1] _099_ VSS VSS VCC VCC _100_ sky130_fd_sc_hd__mux2_1
X_963_ clknet_3_5__leaf_i_clk _022_ VSS VSS VCC VCC o_funct3[0] sky130_fd_sc_hd__dfxtp_2
X_894_ i_pc_next[13] o_pc_next[13] _281_ VSS VSS VCC VCC _407_ sky130_fd_sc_hd__mux2_1
X_946_ clknet_3_4__leaf_i_clk _005_ VSS VSS VCC VCC imm_i\[31\] sky130_fd_sc_hd__dfxtp_1
X_877_ _398_ VSS VSS VCC VCC _044_ sky130_fd_sc_hd__clkbuf_1
X_800_ _353_ VSS VSS VCC VCC _012_ sky130_fd_sc_hd__clkbuf_1
X_731_ i_imm_i[8] imm_i\[8\] _306_ VSS VSS VCC VCC _315_ sky130_fd_sc_hd__mux2_1
X_662_ o_pc[15] i_reg1_data[15] _168_ VSS VSS VCC VCC _271_ sky130_fd_sc_hd__mux2_2
X_593_ imm_i\[7\] i_ret_addr[7] inst_mret VSS VSS VCC VCC _210_ sky130_fd_sc_hd__mux2_1
X_929_ clknet_3_5__leaf_i_clk _085_ VSS VSS VCC VCC imm_i\[14\] sky130_fd_sc_hd__dfxtp_2
X_645_ imm_i\[13\] i_ret_addr[13] _167_ VSS VSS VCC VCC _256_ sky130_fd_sc_hd__mux2_1
X_714_ _281_ VSS VSS VCC VCC _306_ sky130_fd_sc_hd__clkbuf_4
X_576_ _180_ _185_ _191_ _194_ VSS VSS VCC VCC _195_ sky130_fd_sc_hd__o31a_2
X_430_ _108_ VSS VSS VCC VCC o_op1[8] sky130_fd_sc_hd__buf_2
X_628_ o_pc[11] i_reg1_data[11] _168_ VSS VSS VCC VCC _241_ sky130_fd_sc_hd__mux2_2
X_559_ _172_ _178_ _176_ _173_ VSS VSS VCC VCC _180_ sky130_fd_sc_hd__o2bb2a_2
X_413_ op1_sel VSS VSS VCC VCC _099_ sky130_fd_sc_hd__clkbuf_2
X_962_ clknet_3_6__leaf_i_clk _021_ VSS VSS VCC VCC o_reg_write sky130_fd_sc_hd__dfxtp_2
X_893_ _406_ VSS VSS VCC VCC _052_ sky130_fd_sc_hd__clkbuf_1
X_945_ clknet_3_5__leaf_i_clk _004_ VSS VSS VCC VCC imm_i\[30\] sky130_fd_sc_hd__dfxtp_1
X_876_ i_pc_next[4] o_pc_next[4] _390_ VSS VSS VCC VCC _398_ sky130_fd_sc_hd__mux2_1
X_661_ _268_ _270_ VSS VSS VCC VCC o_pc_target[14] sky130_fd_sc_hd__xnor2_4
X_592_ _170_ imm_i\[7\] _208_ VSS VSS VCC VCC _209_ sky130_fd_sc_hd__and3_1
X_730_ _314_ VSS VSS VCC VCC _078_ sky130_fd_sc_hd__clkbuf_1
X_928_ clknet_3_5__leaf_i_clk _084_ VSS VSS VCC VCC imm_i\[13\] sky130_fd_sc_hd__dfxtp_2
X_859_ _388_ VSS VSS VCC VCC _036_ sky130_fd_sc_hd__clkbuf_1
X_644_ imm_i\[13\] VSS VSS VCC VCC _255_ sky130_fd_sc_hd__inv_2
X_575_ _182_ _193_ _190_ VSS VSS VCC VCC _194_ sky130_fd_sc_hd__a21oi_1
X_713_ _305_ VSS VSS VCC VCC _070_ sky130_fd_sc_hd__clkbuf_1
X_627_ _237_ _240_ VSS VSS VCC VCC o_pc_target[10] sky130_fd_sc_hd__xnor2_4
X_558_ _172_ _179_ VSS VSS VCC VCC o_pc_target[2] sky130_fd_sc_hd__xnor2_4
X_489_ _138_ VSS VSS VCC VCC o_op2[5] sky130_fd_sc_hd__buf_2
X_412_ _098_ VSS VSS VCC VCC o_op1[0] sky130_fd_sc_hd__buf_2
X_961_ clknet_3_7__leaf_i_clk _020_ VSS VSS VCC VCC o_res_src[2] sky130_fd_sc_hd__dfxtp_2
X_892_ i_pc_next[12] o_pc_next[12] _281_ VSS VSS VCC VCC _406_ sky130_fd_sc_hd__mux2_1
X_944_ clknet_3_1__leaf_i_clk _003_ VSS VSS VCC VCC imm_i\[29\] sky130_fd_sc_hd__dfxtp_1
X_875_ _397_ VSS VSS VCC VCC _043_ sky130_fd_sc_hd__clkbuf_1
X_660_ _259_ _263_ _269_ VSS VSS VCC VCC _270_ sky130_fd_sc_hd__a21oi_2
X_591_ o_pc[7] i_reg1_data[7] inst_jalr VSS VSS VCC VCC _208_ sky130_fd_sc_hd__mux2_1
X_927_ clknet_3_5__leaf_i_clk _083_ VSS VSS VCC VCC imm_i\[12\] sky130_fd_sc_hd__dfxtp_1
X_858_ i_pc[12] o_pc[12] _379_ VSS VSS VCC VCC _388_ sky130_fd_sc_hd__mux2_1
X_789_ _346_ VSS VSS VCC VCC _008_ sky130_fd_sc_hd__clkbuf_1
X_712_ i_rs2[4] o_rs2[4] _282_ VSS VSS VCC VCC _305_ sky130_fd_sc_hd__mux2_1
X_643_ _253_ _254_ VSS VSS VCC VCC o_pc_target[12] sky130_fd_sc_hd__xnor2_4
X_574_ _186_ _187_ _188_ VSS VSS VCC VCC _193_ sky130_fd_sc_hd__a21o_1
X_626_ _238_ _232_ _239_ VSS VSS VCC VCC _240_ sky130_fd_sc_hd__o21ba_1
X_557_ _173_ _176_ _178_ VSS VSS VCC VCC _179_ sky130_fd_sc_hd__o21ai_2
X_488_ i_reg2_data[5] imm_i\[5\] _132_ VSS VSS VCC VCC _138_ sky130_fd_sc_hd__mux2_1
X_411_ _097_ i_reg1_data[0] VSS VSS VCC VCC _098_ sky130_fd_sc_hd__and2b_1
X_609_ imm_i\[9\] i_ret_addr[9] _167_ VSS VSS VCC VCC _224_ sky130_fd_sc_hd__mux2_1
X_960_ clknet_3_7__leaf_i_clk _019_ VSS VSS VCC VCC o_res_src[1] sky130_fd_sc_hd__dfxtp_2
X_891_ _405_ VSS VSS VCC VCC _051_ sky130_fd_sc_hd__clkbuf_1
X_943_ clknet_3_1__leaf_i_clk _002_ VSS VSS VCC VCC imm_i\[28\] sky130_fd_sc_hd__dfxtp_1
X_874_ i_pc_next[3] o_pc_next[3] _390_ VSS VSS VCC VCC _397_ sky130_fd_sc_hd__mux2_1
X_590_ _206_ _207_ VSS VSS VCC VCC o_pc_target[6] sky130_fd_sc_hd__xnor2_4
X_788_ _289_ _345_ VSS VSS VCC VCC _346_ sky130_fd_sc_hd__and2_1
X_926_ clknet_3_5__leaf_i_clk _082_ VSS VSS VCC VCC imm_i\[11\] sky130_fd_sc_hd__dfxtp_1
X_857_ _387_ VSS VSS VCC VCC _035_ sky130_fd_sc_hd__clkbuf_1
X_642_ _244_ _248_ _242_ VSS VSS VCC VCC _254_ sky130_fd_sc_hd__o21ba_1
X_711_ _304_ VSS VSS VCC VCC _069_ sky130_fd_sc_hd__clkbuf_1
X_573_ _191_ _192_ VSS VSS VCC VCC o_pc_target[4] sky130_fd_sc_hd__xor2_4
X_909_ clknet_3_6__leaf_i_clk _065_ VSS VSS VCC VCC o_rd[4] sky130_fd_sc_hd__dfxtp_2
X_625_ _223_ _227_ VSS VSS VCC VCC _239_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0_i_clk i_clk VSS VSS VCC VCC clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_556_ _170_ _175_ _177_ VSS VSS VCC VCC _178_ sky130_fd_sc_hd__a21o_1
X_487_ _137_ VSS VSS VCC VCC o_op2[4] sky130_fd_sc_hd__buf_2
X_410_ op1_sel VSS VSS VCC VCC _097_ sky130_fd_sc_hd__clkbuf_2
X_608_ imm_i\[9\] VSS VSS VCC VCC _223_ sky130_fd_sc_hd__inv_2
X_539_ _164_ VSS VSS VCC VCC o_op2[29] sky130_fd_sc_hd__buf_2
X_890_ i_pc_next[11] o_pc_next[11] _281_ VSS VSS VCC VCC _405_ sky130_fd_sc_hd__mux2_1
X_942_ clknet_3_1__leaf_i_clk _001_ VSS VSS VCC VCC imm_i\[27\] sky130_fd_sc_hd__dfxtp_1
X_873_ _396_ VSS VSS VCC VCC _042_ sky130_fd_sc_hd__clkbuf_1
X_925_ clknet_3_5__leaf_i_clk _081_ VSS VSS VCC VCC imm_i\[10\] sky130_fd_sc_hd__dfxtp_2
X_787_ i_inst_jal inst_jal _290_ VSS VSS VCC VCC _345_ sky130_fd_sc_hd__mux2_1
X_856_ i_pc[11] o_pc[11] _379_ VSS VSS VCC VCC _387_ sky130_fd_sc_hd__mux2_1
X_641_ _250_ _251_ _252_ VSS VSS VCC VCC _253_ sky130_fd_sc_hd__o21ba_2
X_572_ _180_ _185_ _182_ VSS VSS VCC VCC _192_ sky130_fd_sc_hd__o21ba_1
X_710_ i_rs2[3] o_rs2[3] _282_ VSS VSS VCC VCC _304_ sky130_fd_sc_hd__mux2_1
X_908_ clknet_3_3__leaf_i_clk _064_ VSS VSS VCC VCC o_rd[3] sky130_fd_sc_hd__dfxtp_2
X_839_ i_pc[3] o_pc[3] _339_ VSS VSS VCC VCC _378_ sky130_fd_sc_hd__mux2_1
X_624_ _228_ VSS VSS VCC VCC _238_ sky130_fd_sc_hd__inv_2
X_555_ imm_i\[2\] i_ret_addr[2] inst_mret VSS VSS VCC VCC _177_ sky130_fd_sc_hd__mux2_1
X_486_ i_reg2_data[4] imm_i\[4\] _132_ VSS VSS VCC VCC _137_ sky130_fd_sc_hd__mux2_1
X_607_ _220_ _222_ VSS VSS VCC VCC o_pc_target[8] sky130_fd_sc_hd__xnor2_4
X_538_ i_reg2_data[29] imm_i\[29\] op2_sel VSS VSS VCC VCC _164_ sky130_fd_sc_hd__mux2_1
X_469_ _099_ i_reg1_data[28] VSS VSS VCC VCC _128_ sky130_fd_sc_hd__and2b_1
Xclkbuf_3_2__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_2__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_941_ clknet_3_1__leaf_i_clk _000_ VSS VSS VCC VCC imm_i\[26\] sky130_fd_sc_hd__dfxtp_1
X_872_ i_pc_next[2] o_pc_next[2] _390_ VSS VSS VCC VCC _396_ sky130_fd_sc_hd__mux2_1
X_924_ clknet_3_4__leaf_i_clk _080_ VSS VSS VCC VCC imm_i\[9\] sky130_fd_sc_hd__dfxtp_2
X_786_ _344_ VSS VSS VCC VCC _007_ sky130_fd_sc_hd__clkbuf_1
X_855_ _386_ VSS VSS VCC VCC _034_ sky130_fd_sc_hd__clkbuf_1
X_640_ _225_ imm_i\[12\] _249_ VSS VSS VCC VCC _252_ sky130_fd_sc_hd__and3_1
X_571_ _189_ _190_ VSS VSS VCC VCC _191_ sky130_fd_sc_hd__or2_2
X_838_ _377_ VSS VSS VCC VCC _026_ sky130_fd_sc_hd__clkbuf_1
X_907_ clknet_3_3__leaf_i_clk _063_ VSS VSS VCC VCC o_rd[2] sky130_fd_sc_hd__dfxtp_2
X_769_ i_imm_i[26] imm_i\[26\] _328_ VSS VSS VCC VCC _335_ sky130_fd_sc_hd__mux2_1
X_623_ imm_i\[10\] _234_ _236_ VSS VSS VCC VCC _237_ sky130_fd_sc_hd__a21boi_4
X_554_ _174_ _175_ VSS VSS VCC VCC _176_ sky130_fd_sc_hd__nand2_1
X_485_ _136_ VSS VSS VCC VCC o_op2[3] sky130_fd_sc_hd__buf_2
X_606_ _211_ _215_ _221_ VSS VSS VCC VCC _222_ sky130_fd_sc_hd__o21a_1
X_468_ _127_ VSS VSS VCC VCC o_op1[27] sky130_fd_sc_hd__buf_2
X_537_ _163_ VSS VSS VCC VCC o_op2[28] sky130_fd_sc_hd__buf_2
X_940_ clknet_3_4__leaf_i_clk _096_ VSS VSS VCC VCC imm_i\[25\] sky130_fd_sc_hd__dfxtp_1
X_871_ _395_ VSS VSS VCC VCC _041_ sky130_fd_sc_hd__clkbuf_1
X_923_ clknet_3_4__leaf_i_clk _079_ VSS VSS VCC VCC imm_i\[8\] sky130_fd_sc_hd__dfxtp_1
X_854_ i_pc[10] o_pc[10] _379_ VSS VSS VCC VCC _386_ sky130_fd_sc_hd__mux2_1
X_785_ _289_ _343_ VSS VSS VCC VCC _344_ sky130_fd_sc_hd__and2_1
X_570_ imm_i\[4\] _186_ _187_ VSS VSS VCC VCC _190_ sky130_fd_sc_hd__and3_1
X_768_ _334_ VSS VSS VCC VCC _096_ sky130_fd_sc_hd__clkbuf_1
X_837_ i_pc[2] o_pc[2] _339_ VSS VSS VCC VCC _377_ sky130_fd_sc_hd__mux2_1
X_906_ clknet_3_3__leaf_i_clk _062_ VSS VSS VCC VCC o_rd[1] sky130_fd_sc_hd__dfxtp_2
X_699_ _289_ _297_ VSS VSS VCC VCC _298_ sky130_fd_sc_hd__and2_1
X_622_ _234_ _235_ VSS VSS VCC VCC _236_ sky130_fd_sc_hd__or2_1
X_484_ i_reg2_data[3] imm_i\[3\] _132_ VSS VSS VCC VCC _136_ sky130_fd_sc_hd__mux2_1
X_553_ o_pc[2] i_reg1_data[2] inst_jalr VSS VSS VCC VCC _175_ sky130_fd_sc_hd__mux2_1
X_605_ _209_ VSS VSS VCC VCC _221_ sky130_fd_sc_hd__inv_2
X_467_ _099_ i_reg1_data[27] VSS VSS VCC VCC _127_ sky130_fd_sc_hd__and2b_1
X_536_ i_reg2_data[28] imm_i\[28\] _153_ VSS VSS VCC VCC _163_ sky130_fd_sc_hd__mux2_1
X_519_ _154_ VSS VSS VCC VCC o_op2[19] sky130_fd_sc_hd__buf_2
X_870_ i_pc_next[1] o_pc_next[1] _390_ VSS VSS VCC VCC _395_ sky130_fd_sc_hd__mux2_1
X_784_ i_inst_jalr _168_ _290_ VSS VSS VCC VCC _343_ sky130_fd_sc_hd__mux2_1
X_922_ clknet_3_4__leaf_i_clk _078_ VSS VSS VCC VCC imm_i\[7\] sky130_fd_sc_hd__dfxtp_1
X_853_ _385_ VSS VSS VCC VCC _033_ sky130_fd_sc_hd__clkbuf_1
X_905_ clknet_3_3__leaf_i_clk _061_ VSS VSS VCC VCC o_rd[0] sky130_fd_sc_hd__dfxtp_2
X_767_ i_imm_i[25] imm_i\[25\] _328_ VSS VSS VCC VCC _334_ sky130_fd_sc_hd__mux2_1
X_836_ _376_ VSS VSS VCC VCC _025_ sky130_fd_sc_hd__clkbuf_1
X_698_ i_rd[3] o_rd[3] _290_ VSS VSS VCC VCC _297_ sky130_fd_sc_hd__mux2_1
X_621_ imm_i\[10\] i_ret_addr[10] _167_ VSS VSS VCC VCC _235_ sky130_fd_sc_hd__mux2_1
X_552_ _170_ VSS VSS VCC VCC _174_ sky130_fd_sc_hd__buf_2
X_483_ _135_ VSS VSS VCC VCC o_op2[2] sky130_fd_sc_hd__buf_2
X_819_ _366_ VSS VSS VCC VCC _018_ sky130_fd_sc_hd__clkbuf_1
X_604_ _218_ _219_ VSS VSS VCC VCC _220_ sky130_fd_sc_hd__nor2_2
X_535_ _162_ VSS VSS VCC VCC o_op2[27] sky130_fd_sc_hd__buf_2
X_466_ _126_ VSS VSS VCC VCC o_op1[26] sky130_fd_sc_hd__buf_2
X_518_ i_reg2_data[19] imm_i\[19\] _153_ VSS VSS VCC VCC _154_ sky130_fd_sc_hd__mux2_1
X_449_ _097_ i_reg1_data[18] VSS VSS VCC VCC _118_ sky130_fd_sc_hd__and2b_1
X_921_ clknet_3_1__leaf_i_clk _077_ VSS VSS VCC VCC imm_i\[6\] sky130_fd_sc_hd__dfxtp_2
X_783_ _342_ VSS VSS VCC VCC _006_ sky130_fd_sc_hd__clkbuf_1
X_852_ i_pc[9] o_pc[9] _379_ VSS VSS VCC VCC _385_ sky130_fd_sc_hd__mux2_1
X_904_ clknet_3_2__leaf_i_clk _060_ VSS VSS VCC VCC o_rs1[4] sky130_fd_sc_hd__dfxtp_2
X_766_ _333_ VSS VSS VCC VCC _095_ sky130_fd_sc_hd__clkbuf_1
X_835_ i_pc[1] o_pc[1] _339_ VSS VSS VCC VCC _376_ sky130_fd_sc_hd__mux2_1
X_697_ _296_ VSS VSS VCC VCC _063_ sky130_fd_sc_hd__clkbuf_1
X_551_ imm_i\[2\] VSS VSS VCC VCC _173_ sky130_fd_sc_hd__inv_2
X_620_ _174_ _233_ VSS VSS VCC VCC _234_ sky130_fd_sc_hd__and2_1
Xclkbuf_3_5__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_5__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_482_ i_reg2_data[2] imm_i\[2\] _132_ VSS VSS VCC VCC _135_ sky130_fd_sc_hd__mux2_1
X_818_ _354_ _365_ VSS VSS VCC VCC _366_ sky130_fd_sc_hd__and2_1
X_749_ _324_ VSS VSS VCC VCC _087_ sky130_fd_sc_hd__clkbuf_1
X_603_ _170_ imm_i\[8\] _216_ VSS VSS VCC VCC _219_ sky130_fd_sc_hd__and3_1
X_465_ _099_ i_reg1_data[26] VSS VSS VCC VCC _126_ sky130_fd_sc_hd__and2b_1
X_534_ i_reg2_data[27] imm_i\[27\] _153_ VSS VSS VCC VCC _162_ sky130_fd_sc_hd__mux2_1
X_448_ _117_ VSS VSS VCC VCC o_op1[17] sky130_fd_sc_hd__buf_2
X_517_ op2_sel VSS VSS VCC VCC _153_ sky130_fd_sc_hd__clkbuf_4
X_851_ _384_ VSS VSS VCC VCC _032_ sky130_fd_sc_hd__clkbuf_1
X_920_ clknet_3_1__leaf_i_clk _076_ VSS VSS VCC VCC imm_i\[5\] sky130_fd_sc_hd__dfxtp_1
X_782_ i_op1_src _099_ _339_ VSS VSS VCC VCC _342_ sky130_fd_sc_hd__mux2_1
X_834_ _375_ VSS VSS VCC VCC _024_ sky130_fd_sc_hd__clkbuf_1
X_903_ clknet_3_2__leaf_i_clk _059_ VSS VSS VCC VCC o_rs1[3] sky130_fd_sc_hd__dfxtp_2
X_696_ _289_ _295_ VSS VSS VCC VCC _296_ sky130_fd_sc_hd__and2_1
X_765_ i_imm_i[24] imm_i\[24\] _328_ VSS VSS VCC VCC _333_ sky130_fd_sc_hd__mux2_1
X_550_ _170_ imm_i\[1\] _171_ VSS VSS VCC VCC _172_ sky130_fd_sc_hd__and3_2
X_481_ _134_ VSS VSS VCC VCC o_op2[1] sky130_fd_sc_hd__buf_2
X_817_ i_res_src[0] o_res_src[0] _351_ VSS VSS VCC VCC _365_ sky130_fd_sc_hd__mux2_1
X_748_ i_imm_i[16] imm_i\[16\] _317_ VSS VSS VCC VCC _324_ sky130_fd_sc_hd__mux2_1
X_679_ _284_ VSS VSS VCC VCC _057_ sky130_fd_sc_hd__clkbuf_1
X_602_ _174_ _216_ _217_ VSS VSS VCC VCC _218_ sky130_fd_sc_hd__a21oi_1
X_464_ _125_ VSS VSS VCC VCC o_op1[25] sky130_fd_sc_hd__buf_2
X_533_ _161_ VSS VSS VCC VCC o_op2[26] sky130_fd_sc_hd__buf_2
X_447_ _097_ i_reg1_data[17] VSS VSS VCC VCC _117_ sky130_fd_sc_hd__and2b_1
X_516_ _152_ VSS VSS VCC VCC o_op2[18] sky130_fd_sc_hd__buf_2
X_996_ clknet_3_6__leaf_i_clk _055_ VSS VSS VCC VCC o_pc_next[15] sky130_fd_sc_hd__dfxtp_2
X_781_ _341_ VSS VSS VCC VCC _005_ sky130_fd_sc_hd__clkbuf_1
X_850_ i_pc[8] o_pc[8] _379_ VSS VSS VCC VCC _384_ sky130_fd_sc_hd__mux2_1
X_979_ clknet_3_3__leaf_i_clk _038_ VSS VSS VCC VCC o_pc[14] sky130_fd_sc_hd__dfxtp_2
X_833_ i_funct3[2] o_funct3[2] _339_ VSS VSS VCC VCC _375_ sky130_fd_sc_hd__mux2_1
X_764_ _332_ VSS VSS VCC VCC _094_ sky130_fd_sc_hd__clkbuf_1
X_902_ clknet_3_2__leaf_i_clk _058_ VSS VSS VCC VCC o_rs1[2] sky130_fd_sc_hd__dfxtp_2
X_695_ i_rd[2] o_rd[2] _290_ VSS VSS VCC VCC _295_ sky130_fd_sc_hd__mux2_1
X_480_ i_reg2_data[1] imm_i\[1\] _132_ VSS VSS VCC VCC _134_ sky130_fd_sc_hd__mux2_1
X_816_ _364_ VSS VSS VCC VCC _017_ sky130_fd_sc_hd__clkbuf_1
X_747_ _323_ VSS VSS VCC VCC _086_ sky130_fd_sc_hd__clkbuf_1
X_678_ i_rs1[1] o_rs1[1] _282_ VSS VSS VCC VCC _284_ sky130_fd_sc_hd__mux2_1
X_601_ imm_i\[8\] i_ret_addr[8] inst_mret VSS VSS VCC VCC _217_ sky130_fd_sc_hd__mux2_1
X_463_ _099_ i_reg1_data[25] VSS VSS VCC VCC _125_ sky130_fd_sc_hd__and2b_1
X_532_ i_reg2_data[26] imm_i\[26\] _153_ VSS VSS VCC VCC _161_ sky130_fd_sc_hd__mux2_1
X_515_ i_reg2_data[18] imm_i\[18\] _142_ VSS VSS VCC VCC _152_ sky130_fd_sc_hd__mux2_1
X_446_ _116_ VSS VSS VCC VCC o_op1[16] sky130_fd_sc_hd__buf_2
X_995_ clknet_3_6__leaf_i_clk _054_ VSS VSS VCC VCC o_pc_next[14] sky130_fd_sc_hd__dfxtp_2
X_429_ i_reg1_data[8] o_pc[8] _102_ VSS VSS VCC VCC _108_ sky130_fd_sc_hd__mux2_1
X_780_ i_imm_i[31] imm_i\[31\] _339_ VSS VSS VCC VCC _341_ sky130_fd_sc_hd__mux2_1
X_978_ clknet_3_3__leaf_i_clk _037_ VSS VSS VCC VCC o_pc[13] sky130_fd_sc_hd__dfxtp_2
X_901_ clknet_3_2__leaf_i_clk _057_ VSS VSS VCC VCC o_rs1[1] sky130_fd_sc_hd__dfxtp_2
X_832_ _374_ VSS VSS VCC VCC _023_ sky130_fd_sc_hd__clkbuf_1
X_763_ i_imm_i[23] imm_i\[23\] _328_ VSS VSS VCC VCC _332_ sky130_fd_sc_hd__mux2_1
X_694_ _294_ VSS VSS VCC VCC _062_ sky130_fd_sc_hd__clkbuf_1
X_815_ _354_ _363_ VSS VSS VCC VCC _364_ sky130_fd_sc_hd__and2_1
X_746_ i_imm_i[15] imm_i\[15\] _317_ VSS VSS VCC VCC _323_ sky130_fd_sc_hd__mux2_1
X_677_ _283_ VSS VSS VCC VCC _056_ sky130_fd_sc_hd__clkbuf_1
X_531_ _160_ VSS VSS VCC VCC o_op2[25] sky130_fd_sc_hd__buf_2
X_600_ o_pc[8] i_reg1_data[8] inst_jalr VSS VSS VCC VCC _216_ sky130_fd_sc_hd__mux2_1
X_462_ _124_ VSS VSS VCC VCC o_op1[24] sky130_fd_sc_hd__buf_2
X_729_ i_imm_i[7] imm_i\[7\] _306_ VSS VSS VCC VCC _314_ sky130_fd_sc_hd__mux2_1
X_514_ _151_ VSS VSS VCC VCC o_op2[17] sky130_fd_sc_hd__buf_2
X_445_ _097_ i_reg1_data[16] VSS VSS VCC VCC _116_ sky130_fd_sc_hd__and2b_1
X_994_ clknet_3_6__leaf_i_clk _053_ VSS VSS VCC VCC o_pc_next[13] sky130_fd_sc_hd__dfxtp_2
X_428_ _107_ VSS VSS VCC VCC o_op1[7] sky130_fd_sc_hd__buf_2
X_977_ clknet_3_2__leaf_i_clk _036_ VSS VSS VCC VCC o_pc[12] sky130_fd_sc_hd__dfxtp_2
X_831_ i_funct3[1] o_funct3[1] _339_ VSS VSS VCC VCC _374_ sky130_fd_sc_hd__mux2_1
X_900_ clknet_3_2__leaf_i_clk _056_ VSS VSS VCC VCC o_rs1[0] sky130_fd_sc_hd__dfxtp_2
X_693_ _289_ _293_ VSS VSS VCC VCC _294_ sky130_fd_sc_hd__and2_1
X_762_ _331_ VSS VSS VCC VCC _093_ sky130_fd_sc_hd__clkbuf_1
X_814_ i_inst_store o_store _351_ VSS VSS VCC VCC _363_ sky130_fd_sc_hd__mux2_1
X_745_ _322_ VSS VSS VCC VCC _085_ sky130_fd_sc_hd__clkbuf_1
X_676_ i_rs1[0] o_rs1[0] _282_ VSS VSS VCC VCC _283_ sky130_fd_sc_hd__mux2_1
X_461_ _097_ i_reg1_data[24] VSS VSS VCC VCC _124_ sky130_fd_sc_hd__and2b_1
X_530_ i_reg2_data[25] imm_i\[25\] _153_ VSS VSS VCC VCC _160_ sky130_fd_sc_hd__mux2_1
X_659_ _255_ _258_ VSS VSS VCC VCC _269_ sky130_fd_sc_hd__nor2_1
X_728_ _313_ VSS VSS VCC VCC _077_ sky130_fd_sc_hd__clkbuf_1
X_444_ _115_ VSS VSS VCC VCC o_op1[15] sky130_fd_sc_hd__buf_2
X_513_ i_reg2_data[17] imm_i\[17\] _142_ VSS VSS VCC VCC _151_ sky130_fd_sc_hd__mux2_1
X_993_ clknet_3_6__leaf_i_clk _052_ VSS VSS VCC VCC o_pc_next[12] sky130_fd_sc_hd__dfxtp_2
X_427_ i_reg1_data[7] o_pc[7] _102_ VSS VSS VCC VCC _107_ sky130_fd_sc_hd__mux2_1
X_976_ clknet_3_2__leaf_i_clk _035_ VSS VSS VCC VCC o_pc[11] sky130_fd_sc_hd__dfxtp_2
X_830_ _373_ VSS VSS VCC VCC _022_ sky130_fd_sc_hd__clkbuf_1
X_761_ i_imm_i[22] imm_i\[22\] _328_ VSS VSS VCC VCC _331_ sky130_fd_sc_hd__mux2_1
X_692_ i_rd[1] o_rd[1] _290_ VSS VSS VCC VCC _293_ sky130_fd_sc_hd__mux2_1
X_959_ clknet_3_6__leaf_i_clk _018_ VSS VSS VCC VCC o_res_src[0] sky130_fd_sc_hd__dfxtp_2
X_813_ _362_ VSS VSS VCC VCC _016_ sky130_fd_sc_hd__clkbuf_1
X_744_ i_imm_i[14] imm_i\[14\] _317_ VSS VSS VCC VCC _322_ sky130_fd_sc_hd__mux2_1
X_675_ _281_ VSS VSS VCC VCC _282_ sky130_fd_sc_hd__clkbuf_4
X_460_ _123_ VSS VSS VCC VCC o_op1[23] sky130_fd_sc_hd__buf_2
X_727_ i_imm_i[6] imm_i\[6\] _306_ VSS VSS VCC VCC _313_ sky130_fd_sc_hd__mux2_1
X_658_ _266_ _267_ VSS VSS VCC VCC _268_ sky130_fd_sc_hd__nor2_2
X_589_ _195_ _199_ _197_ VSS VSS VCC VCC _207_ sky130_fd_sc_hd__o21ba_1
X_443_ i_reg1_data[15] o_pc[15] op1_sel VSS VSS VCC VCC _115_ sky130_fd_sc_hd__mux2_1
X_512_ _150_ VSS VSS VCC VCC o_op2[16] sky130_fd_sc_hd__buf_2
X_992_ clknet_3_6__leaf_i_clk _051_ VSS VSS VCC VCC o_pc_next[11] sky130_fd_sc_hd__dfxtp_2
X_426_ _106_ VSS VSS VCC VCC o_op1[6] sky130_fd_sc_hd__buf_2
X_975_ clknet_3_2__leaf_i_clk _034_ VSS VSS VCC VCC o_pc[10] sky130_fd_sc_hd__dfxtp_2
X_760_ _330_ VSS VSS VCC VCC _092_ sky130_fd_sc_hd__clkbuf_1
X_691_ _292_ VSS VSS VCC VCC _061_ sky130_fd_sc_hd__clkbuf_1
X_958_ clknet_3_7__leaf_i_clk _017_ VSS VSS VCC VCC o_store sky130_fd_sc_hd__dfxtp_2
X_889_ _404_ VSS VSS VCC VCC _050_ sky130_fd_sc_hd__clkbuf_1
X_812_ _354_ _361_ VSS VSS VCC VCC _362_ sky130_fd_sc_hd__and2_1
X_743_ _321_ VSS VSS VCC VCC _084_ sky130_fd_sc_hd__clkbuf_1
X_674_ _280_ VSS VSS VCC VCC _281_ sky130_fd_sc_hd__clkbuf_4
X_657_ _225_ imm_i\[14\] _264_ VSS VSS VCC VCC _267_ sky130_fd_sc_hd__and3_1
X_726_ _312_ VSS VSS VCC VCC _076_ sky130_fd_sc_hd__clkbuf_1
X_588_ imm_i\[6\] _203_ _205_ VSS VSS VCC VCC _206_ sky130_fd_sc_hd__a21boi_4
X_511_ i_reg2_data[16] imm_i\[16\] _142_ VSS VSS VCC VCC _150_ sky130_fd_sc_hd__mux2_1
X_442_ _114_ VSS VSS VCC VCC o_op1[14] sky130_fd_sc_hd__buf_2
X_709_ _303_ VSS VSS VCC VCC _068_ sky130_fd_sc_hd__clkbuf_1
X_991_ clknet_3_3__leaf_i_clk _050_ VSS VSS VCC VCC o_pc_next[10] sky130_fd_sc_hd__dfxtp_2
X_425_ i_reg1_data[6] o_pc[6] _102_ VSS VSS VCC VCC _106_ sky130_fd_sc_hd__mux2_1
X_974_ clknet_3_2__leaf_i_clk _033_ VSS VSS VCC VCC o_pc[9] sky130_fd_sc_hd__dfxtp_2
X_690_ _289_ _291_ VSS VSS VCC VCC _292_ sky130_fd_sc_hd__and2_1
X_957_ clknet_3_7__leaf_i_clk _016_ VSS VSS VCC VCC o_alu_ctrl[4] sky130_fd_sc_hd__dfxtp_2
X_888_ i_pc_next[10] o_pc_next[10] _281_ VSS VSS VCC VCC _404_ sky130_fd_sc_hd__mux2_1
X_811_ i_alu_ctrl[4] o_alu_ctrl[4] _351_ VSS VSS VCC VCC _361_ sky130_fd_sc_hd__mux2_1
X_742_ i_imm_i[13] imm_i\[13\] _317_ VSS VSS VCC VCC _321_ sky130_fd_sc_hd__mux2_1
X_673_ _279_ VSS VSS VCC VCC _280_ sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_3_1__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_1__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_656_ _225_ _264_ _265_ VSS VSS VCC VCC _266_ sky130_fd_sc_hd__a21oi_1
X_725_ i_imm_i[5] imm_i\[5\] _306_ VSS VSS VCC VCC _312_ sky130_fd_sc_hd__mux2_1
X_587_ _174_ _201_ _202_ _204_ VSS VSS VCC VCC _205_ sky130_fd_sc_hd__a31o_1
X_441_ i_reg1_data[14] o_pc[14] op1_sel VSS VSS VCC VCC _114_ sky130_fd_sc_hd__mux2_1
X_510_ _149_ VSS VSS VCC VCC o_op2[15] sky130_fd_sc_hd__buf_2
X_639_ imm_i\[12\] i_ret_addr[12] _167_ VSS VSS VCC VCC _251_ sky130_fd_sc_hd__mux2_1
X_708_ i_rs2[2] o_rs2[2] _282_ VSS VSS VCC VCC _303_ sky130_fd_sc_hd__mux2_1
X_990_ clknet_3_3__leaf_i_clk _049_ VSS VSS VCC VCC o_pc_next[9] sky130_fd_sc_hd__dfxtp_2
X_424_ _105_ VSS VSS VCC VCC o_op1[5] sky130_fd_sc_hd__buf_2
X_973_ clknet_3_0__leaf_i_clk _032_ VSS VSS VCC VCC o_pc[8] sky130_fd_sc_hd__dfxtp_2
X_956_ clknet_3_7__leaf_i_clk _015_ VSS VSS VCC VCC o_alu_ctrl[3] sky130_fd_sc_hd__dfxtp_2
X_887_ _403_ VSS VSS VCC VCC _049_ sky130_fd_sc_hd__clkbuf_1
X_810_ _360_ VSS VSS VCC VCC _015_ sky130_fd_sc_hd__clkbuf_1
X_672_ i_stall i_flush i_reset_n VSS VSS VCC VCC _279_ sky130_fd_sc_hd__or3b_1
X_741_ _320_ VSS VSS VCC VCC _083_ sky130_fd_sc_hd__clkbuf_1
X_939_ clknet_3_0__leaf_i_clk _095_ VSS VSS VCC VCC imm_i\[24\] sky130_fd_sc_hd__dfxtp_1
X_724_ _311_ VSS VSS VCC VCC _075_ sky130_fd_sc_hd__clkbuf_1
X_655_ imm_i\[14\] i_ret_addr[14] _167_ VSS VSS VCC VCC _265_ sky130_fd_sc_hd__mux2_1
X_586_ imm_i\[6\] i_ret_addr[6] inst_mret VSS VSS VCC VCC _204_ sky130_fd_sc_hd__mux2_1
X_440_ _113_ VSS VSS VCC VCC o_op1[13] sky130_fd_sc_hd__buf_2
X_707_ _302_ VSS VSS VCC VCC _067_ sky130_fd_sc_hd__clkbuf_1
X_638_ _225_ _249_ VSS VSS VCC VCC _250_ sky130_fd_sc_hd__and2_1
X_569_ _186_ _187_ _188_ VSS VSS VCC VCC _189_ sky130_fd_sc_hd__a21oi_1
X_423_ i_reg1_data[5] o_pc[5] _102_ VSS VSS VCC VCC _105_ sky130_fd_sc_hd__mux2_1
X_972_ clknet_3_0__leaf_i_clk _031_ VSS VSS VCC VCC o_pc[7] sky130_fd_sc_hd__dfxtp_2
X_955_ clknet_3_7__leaf_i_clk _014_ VSS VSS VCC VCC o_alu_ctrl[2] sky130_fd_sc_hd__dfxtp_2
X_886_ i_pc_next[9] o_pc_next[9] _281_ VSS VSS VCC VCC _403_ sky130_fd_sc_hd__mux2_1
X_740_ i_imm_i[12] imm_i\[12\] _317_ VSS VSS VCC VCC _320_ sky130_fd_sc_hd__mux2_1
X_671_ _172_ _278_ VSS VSS VCC VCC o_pc_target[1] sky130_fd_sc_hd__nor2_4
X_869_ _394_ VSS VSS VCC VCC _040_ sky130_fd_sc_hd__clkbuf_1
X_938_ clknet_3_0__leaf_i_clk _094_ VSS VSS VCC VCC imm_i\[23\] sky130_fd_sc_hd__dfxtp_1
X_723_ i_imm_i[4] imm_i\[4\] _306_ VSS VSS VCC VCC _311_ sky130_fd_sc_hd__mux2_1
X_654_ o_pc[14] i_reg1_data[14] _168_ VSS VSS VCC VCC _264_ sky130_fd_sc_hd__mux2_2
X_585_ _174_ _201_ _202_ VSS VSS VCC VCC _203_ sky130_fd_sc_hd__and3_1
X_637_ o_pc[12] i_reg1_data[12] _168_ VSS VSS VCC VCC _249_ sky130_fd_sc_hd__mux2_1
X_706_ i_rs2[1] o_rs2[1] _282_ VSS VSS VCC VCC _302_ sky130_fd_sc_hd__mux2_1
X_568_ imm_i\[4\] i_ret_addr[4] inst_mret VSS VSS VCC VCC _188_ sky130_fd_sc_hd__mux2_1
X_499_ i_reg2_data[10] imm_i\[10\] _142_ VSS VSS VCC VCC _144_ sky130_fd_sc_hd__mux2_1
X_422_ _104_ VSS VSS VCC VCC o_op1[4] sky130_fd_sc_hd__buf_2
X_971_ clknet_3_0__leaf_i_clk _030_ VSS VSS VCC VCC o_pc[6] sky130_fd_sc_hd__dfxtp_2
X_954_ clknet_3_7__leaf_i_clk _013_ VSS VSS VCC VCC o_alu_ctrl[1] sky130_fd_sc_hd__dfxtp_2
X_885_ _402_ VSS VSS VCC VCC _048_ sky130_fd_sc_hd__clkbuf_1
X_670_ _225_ _171_ _277_ VSS VSS VCC VCC _278_ sky130_fd_sc_hd__a21oi_1
X_868_ _354_ _393_ VSS VSS VCC VCC _394_ sky130_fd_sc_hd__and2_1
X_799_ _289_ _352_ VSS VSS VCC VCC _353_ sky130_fd_sc_hd__and2_1
X_937_ clknet_3_0__leaf_i_clk _093_ VSS VSS VCC VCC imm_i\[22\] sky130_fd_sc_hd__dfxtp_1
X_653_ _259_ _263_ VSS VSS VCC VCC o_pc_target[13] sky130_fd_sc_hd__xor2_4
X_722_ _310_ VSS VSS VCC VCC _074_ sky130_fd_sc_hd__clkbuf_1
X_584_ inst_jalr o_pc[6] VSS VSS VCC VCC _202_ sky130_fd_sc_hd__or2_1
X_636_ _245_ _248_ VSS VSS VCC VCC o_pc_target[11] sky130_fd_sc_hd__xnor2_4
X_567_ inst_jalr o_pc[4] inst_mret VSS VSS VCC VCC _187_ sky130_fd_sc_hd__o21ba_1
X_705_ _301_ VSS VSS VCC VCC _066_ sky130_fd_sc_hd__clkbuf_1
X_498_ _143_ VSS VSS VCC VCC o_op2[9] sky130_fd_sc_hd__buf_2
X_421_ i_reg1_data[4] o_pc[4] _102_ VSS VSS VCC VCC _104_ sky130_fd_sc_hd__mux2_1
X_619_ o_pc[10] i_reg1_data[10] _168_ VSS VSS VCC VCC _233_ sky130_fd_sc_hd__mux2_1
X_970_ clknet_3_0__leaf_i_clk _029_ VSS VSS VCC VCC o_pc[5] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_3_4__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_4__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_953_ clknet_3_7__leaf_i_clk _012_ VSS VSS VCC VCC o_alu_ctrl[0] sky130_fd_sc_hd__dfxtp_2
X_884_ i_pc_next[8] o_pc_next[8] _390_ VSS VSS VCC VCC _402_ sky130_fd_sc_hd__mux2_1
X_936_ clknet_3_0__leaf_i_clk _092_ VSS VSS VCC VCC imm_i\[21\] sky130_fd_sc_hd__dfxtp_1
X_867_ i_to_trap o_to_trap i_stall VSS VSS VCC VCC _393_ sky130_fd_sc_hd__mux2_1
X_798_ i_alu_ctrl[0] o_alu_ctrl[0] _351_ VSS VSS VCC VCC _352_ sky130_fd_sc_hd__mux2_1
X_652_ _232_ _246_ _260_ _262_ VSS VSS VCC VCC _263_ sky130_fd_sc_hd__o31ai_4
X_721_ i_imm_i[3] imm_i\[3\] _306_ VSS VSS VCC VCC _310_ sky130_fd_sc_hd__mux2_1
X_583_ i_reg1_data[6] _168_ VSS VSS VCC VCC _201_ sky130_fd_sc_hd__or2b_1
X_919_ clknet_3_1__leaf_i_clk _075_ VSS VSS VCC VCC imm_i\[4\] sky130_fd_sc_hd__dfxtp_1
X_704_ i_rs2[0] o_rs2[0] _282_ VSS VSS VCC VCC _301_ sky130_fd_sc_hd__mux2_1
X_635_ _232_ _246_ _247_ VSS VSS VCC VCC _248_ sky130_fd_sc_hd__o21ba_2
X_566_ i_reg1_data[4] inst_jalr VSS VSS VCC VCC _186_ sky130_fd_sc_hd__or2b_1
X_497_ i_reg2_data[9] imm_i\[9\] _142_ VSS VSS VCC VCC _143_ sky130_fd_sc_hd__mux2_1
X_420_ _103_ VSS VSS VCC VCC o_op1[3] sky130_fd_sc_hd__buf_2
X_618_ _228_ _232_ VSS VSS VCC VCC o_pc_target[9] sky130_fd_sc_hd__xnor2_4
X_549_ o_pc[1] i_reg1_data[1] inst_jalr VSS VSS VCC VCC _171_ sky130_fd_sc_hd__mux2_1
X_883_ _401_ VSS VSS VCC VCC _047_ sky130_fd_sc_hd__clkbuf_1
X_952_ clknet_3_0__leaf_i_clk _011_ VSS VSS VCC VCC op2_sel sky130_fd_sc_hd__dfxtp_1
X_935_ clknet_3_0__leaf_i_clk _091_ VSS VSS VCC VCC imm_i\[20\] sky130_fd_sc_hd__dfxtp_1
X_866_ _392_ VSS VSS VCC VCC _039_ sky130_fd_sc_hd__clkbuf_1
X_797_ i_stall VSS VSS VCC VCC _351_ sky130_fd_sc_hd__clkbuf_4
X_720_ _309_ VSS VSS VCC VCC _073_ sky130_fd_sc_hd__clkbuf_1
X_651_ _245_ _247_ _253_ _261_ _252_ VSS VSS VCC VCC _262_ sky130_fd_sc_hd__a311oi_4
X_582_ _195_ _200_ VSS VSS VCC VCC o_pc_target[5] sky130_fd_sc_hd__xnor2_4
X_918_ clknet_3_4__leaf_i_clk _074_ VSS VSS VCC VCC imm_i\[3\] sky130_fd_sc_hd__dfxtp_1
X_849_ _383_ VSS VSS VCC VCC _031_ sky130_fd_sc_hd__clkbuf_1
X_634_ imm_i\[10\] _234_ _236_ _239_ VSS VSS VCC VCC _247_ sky130_fd_sc_hd__a22o_1
X_703_ _300_ VSS VSS VCC VCC _065_ sky130_fd_sc_hd__clkbuf_1
X_565_ _180_ _185_ VSS VSS VCC VCC o_pc_target[3] sky130_fd_sc_hd__xor2_4
X_496_ op2_sel VSS VSS VCC VCC _142_ sky130_fd_sc_hd__clkbuf_4
X_617_ _195_ _213_ _229_ _231_ VSS VSS VCC VCC _232_ sky130_fd_sc_hd__o31a_4
X_548_ inst_mret VSS VSS VCC VCC _170_ sky130_fd_sc_hd__inv_2
X_479_ _133_ VSS VSS VCC VCC o_op2[0] sky130_fd_sc_hd__buf_2
X_951_ clknet_3_5__leaf_i_clk _010_ VSS VSS VCC VCC inst_mret sky130_fd_sc_hd__dfxtp_4
X_882_ i_pc_next[7] o_pc_next[7] _390_ VSS VSS VCC VCC _401_ sky130_fd_sc_hd__mux2_1
X_934_ clknet_3_4__leaf_i_clk _090_ VSS VSS VCC VCC imm_i\[19\] sky130_fd_sc_hd__dfxtp_1
X_796_ _350_ VSS VSS VCC VCC _011_ sky130_fd_sc_hd__clkbuf_1
X_865_ i_pc[15] o_pc[15] _390_ VSS VSS VCC VCC _392_ sky130_fd_sc_hd__mux2_1
X_650_ _250_ _251_ _242_ VSS VSS VCC VCC _261_ sky130_fd_sc_hd__o21a_1
X_581_ _197_ _199_ VSS VSS VCC VCC _200_ sky130_fd_sc_hd__nor2_2
X_779_ _340_ VSS VSS VCC VCC _004_ sky130_fd_sc_hd__clkbuf_1
X_917_ clknet_3_4__leaf_i_clk _073_ VSS VSS VCC VCC imm_i\[2\] sky130_fd_sc_hd__dfxtp_2
X_848_ i_pc[7] o_pc[7] _379_ VSS VSS VCC VCC _383_ sky130_fd_sc_hd__mux2_1
X_633_ _228_ _237_ VSS VSS VCC VCC _246_ sky130_fd_sc_hd__nand2_1
X_702_ _289_ _299_ VSS VSS VCC VCC _300_ sky130_fd_sc_hd__and2_1
X_564_ _182_ _184_ VSS VSS VCC VCC _185_ sky130_fd_sc_hd__or2_2
X_495_ _141_ VSS VSS VCC VCC o_op2[8] sky130_fd_sc_hd__buf_2
X_547_ _169_ VSS VSS VCC VCC o_inst_jal_jalr sky130_fd_sc_hd__buf_2
X_616_ _221_ _218_ _229_ _214_ _230_ VSS VSS VCC VCC _231_ sky130_fd_sc_hd__o221a_1
X_478_ i_reg2_data[0] imm_i\[0\] _132_ VSS VSS VCC VCC _133_ sky130_fd_sc_hd__mux2_1
X_950_ clknet_3_7__leaf_i_clk _009_ VSS VSS VCC VCC o_inst_branch sky130_fd_sc_hd__dfxtp_2
X_881_ _400_ VSS VSS VCC VCC _046_ sky130_fd_sc_hd__clkbuf_1
X_933_ clknet_3_4__leaf_i_clk _089_ VSS VSS VCC VCC imm_i\[18\] sky130_fd_sc_hd__dfxtp_1
X_795_ i_op2_src _132_ _339_ VSS VSS VCC VCC _350_ sky130_fd_sc_hd__mux2_1
X_864_ _391_ VSS VSS VCC VCC _038_ sky130_fd_sc_hd__clkbuf_1
X_580_ _174_ _196_ _198_ VSS VSS VCC VCC _199_ sky130_fd_sc_hd__a21oi_1
X_916_ clknet_3_1__leaf_i_clk _072_ VSS VSS VCC VCC imm_i\[1\] sky130_fd_sc_hd__dfxtp_1
X_778_ i_imm_i[30] imm_i\[30\] _339_ VSS VSS VCC VCC _340_ sky130_fd_sc_hd__mux2_1
X_847_ _382_ VSS VSS VCC VCC _030_ sky130_fd_sc_hd__clkbuf_1
X_632_ _242_ _244_ VSS VSS VCC VCC _245_ sky130_fd_sc_hd__nor2_4
X_701_ i_rd[4] o_rd[4] _290_ VSS VSS VCC VCC _299_ sky130_fd_sc_hd__mux2_1
X_563_ _174_ _181_ _183_ VSS VSS VCC VCC _184_ sky130_fd_sc_hd__a21oi_1
X_494_ i_reg2_data[8] imm_i\[8\] _132_ VSS VSS VCC VCC _141_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_7__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_7__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_546_ _167_ inst_jal _168_ VSS VSS VCC VCC _169_ sky130_fd_sc_hd__or3_1
X_615_ _219_ VSS VSS VCC VCC _230_ sky130_fd_sc_hd__inv_2
X_477_ op2_sel VSS VSS VCC VCC _132_ sky130_fd_sc_hd__clkbuf_4
X_529_ _159_ VSS VSS VCC VCC o_op2[24] sky130_fd_sc_hd__buf_2
X_880_ i_pc_next[6] o_pc_next[6] _390_ VSS VSS VCC VCC _400_ sky130_fd_sc_hd__mux2_1
X_932_ clknet_3_4__leaf_i_clk _088_ VSS VSS VCC VCC imm_i\[17\] sky130_fd_sc_hd__dfxtp_1
X_863_ i_pc[14] o_pc[14] _390_ VSS VSS VCC VCC _391_ sky130_fd_sc_hd__mux2_1
X_794_ _290_ _225_ _349_ VSS VSS VCC VCC _010_ sky130_fd_sc_hd__a21oi_1
X_915_ clknet_3_1__leaf_i_clk _071_ VSS VSS VCC VCC imm_i\[0\] sky130_fd_sc_hd__dfxtp_1
X_846_ i_pc[6] o_pc[6] _379_ VSS VSS VCC VCC _382_ sky130_fd_sc_hd__mux2_1
X_777_ _280_ VSS VSS VCC VCC _339_ sky130_fd_sc_hd__buf_4
X_700_ _298_ VSS VSS VCC VCC _064_ sky130_fd_sc_hd__clkbuf_1
X_631_ _225_ _241_ _243_ VSS VSS VCC VCC _244_ sky130_fd_sc_hd__a21oi_2
X_562_ imm_i\[3\] i_ret_addr[3] inst_mret VSS VSS VCC VCC _183_ sky130_fd_sc_hd__mux2_1
X_493_ _140_ VSS VSS VCC VCC o_op2[7] sky130_fd_sc_hd__buf_2
X_829_ i_funct3[0] o_funct3[0] _339_ VSS VSS VCC VCC _373_ sky130_fd_sc_hd__mux2_1
X_614_ _209_ _211_ _218_ _219_ VSS VSS VCC VCC _229_ sky130_fd_sc_hd__or4_1
X_476_ _131_ VSS VSS VCC VCC o_op1[31] sky130_fd_sc_hd__buf_2
X_545_ inst_jalr VSS VSS VCC VCC _168_ sky130_fd_sc_hd__buf_4
X_459_ _097_ i_reg1_data[23] VSS VSS VCC VCC _123_ sky130_fd_sc_hd__and2b_1
X_528_ i_reg2_data[24] imm_i\[24\] _153_ VSS VSS VCC VCC _159_ sky130_fd_sc_hd__mux2_1
X_931_ clknet_3_4__leaf_i_clk _087_ VSS VSS VCC VCC imm_i\[16\] sky130_fd_sc_hd__dfxtp_1
X_862_ _280_ VSS VSS VCC VCC _390_ sky130_fd_sc_hd__clkbuf_4
X_793_ _290_ i_inst_mret _289_ VSS VSS VCC VCC _349_ sky130_fd_sc_hd__o21ai_1
X_845_ _381_ VSS VSS VCC VCC _029_ sky130_fd_sc_hd__clkbuf_1
X_914_ clknet_3_3__leaf_i_clk _070_ VSS VSS VCC VCC o_rs2[4] sky130_fd_sc_hd__dfxtp_2
X_776_ _338_ VSS VSS VCC VCC _003_ sky130_fd_sc_hd__clkbuf_1
X_630_ imm_i\[11\] i_ret_addr[11] _167_ VSS VSS VCC VCC _243_ sky130_fd_sc_hd__mux2_1
X_561_ _170_ imm_i\[3\] _181_ VSS VSS VCC VCC _182_ sky130_fd_sc_hd__and3_1
X_492_ i_reg2_data[7] imm_i\[7\] _132_ VSS VSS VCC VCC _140_ sky130_fd_sc_hd__mux2_1
X_828_ _372_ VSS VSS VCC VCC _021_ sky130_fd_sc_hd__clkbuf_1
X_759_ i_imm_i[21] imm_i\[21\] _328_ VSS VSS VCC VCC _330_ sky130_fd_sc_hd__mux2_1
X_613_ _223_ _224_ _227_ VSS VSS VCC VCC _228_ sky130_fd_sc_hd__mux2_2
X_544_ inst_mret VSS VSS VCC VCC _167_ sky130_fd_sc_hd__clkbuf_4
X_475_ _099_ i_reg1_data[31] VSS VSS VCC VCC _131_ sky130_fd_sc_hd__and2b_1
X_527_ _158_ VSS VSS VCC VCC o_op2[23] sky130_fd_sc_hd__buf_2
X_458_ _122_ VSS VSS VCC VCC o_op1[22] sky130_fd_sc_hd__buf_2
X_930_ clknet_3_5__leaf_i_clk _086_ VSS VSS VCC VCC imm_i\[15\] sky130_fd_sc_hd__dfxtp_2
X_792_ _348_ VSS VSS VCC VCC _009_ sky130_fd_sc_hd__clkbuf_1
X_861_ _389_ VSS VSS VCC VCC _037_ sky130_fd_sc_hd__clkbuf_1
X_913_ clknet_3_3__leaf_i_clk _069_ VSS VSS VCC VCC o_rs2[3] sky130_fd_sc_hd__dfxtp_2
X_844_ i_pc[5] o_pc[5] _379_ VSS VSS VCC VCC _381_ sky130_fd_sc_hd__mux2_1
X_775_ i_imm_i[29] imm_i\[29\] _328_ VSS VSS VCC VCC _338_ sky130_fd_sc_hd__mux2_1
X_560_ o_pc[3] i_reg1_data[3] inst_jalr VSS VSS VCC VCC _181_ sky130_fd_sc_hd__mux2_1
X_491_ _139_ VSS VSS VCC VCC o_op2[6] sky130_fd_sc_hd__buf_2
X_827_ _354_ _371_ VSS VSS VCC VCC _372_ sky130_fd_sc_hd__and2_1
X_689_ i_rd[0] o_rd[0] _290_ VSS VSS VCC VCC _291_ sky130_fd_sc_hd__mux2_1
X_758_ _329_ VSS VSS VCC VCC _091_ sky130_fd_sc_hd__clkbuf_1
X_612_ _225_ _226_ VSS VSS VCC VCC _227_ sky130_fd_sc_hd__nand2_1
X_543_ _166_ VSS VSS VCC VCC o_op2[31] sky130_fd_sc_hd__buf_2
X_474_ _130_ VSS VSS VCC VCC o_op1[30] sky130_fd_sc_hd__buf_2
X_526_ i_reg2_data[23] imm_i\[23\] _153_ VSS VSS VCC VCC _158_ sky130_fd_sc_hd__mux2_1
X_457_ _097_ i_reg1_data[22] VSS VSS VCC VCC _122_ sky130_fd_sc_hd__and2b_1
Xclkbuf_3_0__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_0__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_509_ i_reg2_data[15] imm_i\[15\] _142_ VSS VSS VCC VCC _149_ sky130_fd_sc_hd__mux2_1
X_791_ _289_ _347_ VSS VSS VCC VCC _348_ sky130_fd_sc_hd__and2_1
X_860_ i_pc[13] o_pc[13] _379_ VSS VSS VCC VCC _389_ sky130_fd_sc_hd__mux2_1
X_989_ clknet_3_6__leaf_i_clk _048_ VSS VSS VCC VCC o_pc_next[8] sky130_fd_sc_hd__dfxtp_2
X_843_ _380_ VSS VSS VCC VCC _028_ sky130_fd_sc_hd__clkbuf_1
X_912_ clknet_3_2__leaf_i_clk _068_ VSS VSS VCC VCC o_rs2[2] sky130_fd_sc_hd__dfxtp_2
X_774_ _337_ VSS VSS VCC VCC _002_ sky130_fd_sc_hd__clkbuf_1
X_490_ i_reg2_data[6] imm_i\[6\] _132_ VSS VSS VCC VCC _139_ sky130_fd_sc_hd__mux2_1
X_826_ i_reg_write o_reg_write _351_ VSS VSS VCC VCC _371_ sky130_fd_sc_hd__mux2_1
X_688_ i_stall VSS VSS VCC VCC _290_ sky130_fd_sc_hd__clkbuf_4
X_757_ i_imm_i[20] imm_i\[20\] _328_ VSS VSS VCC VCC _329_ sky130_fd_sc_hd__mux2_1
X_473_ _099_ i_reg1_data[30] VSS VSS VCC VCC _130_ sky130_fd_sc_hd__and2b_1
X_611_ o_pc[9] i_reg1_data[9] _168_ VSS VSS VCC VCC _226_ sky130_fd_sc_hd__mux2_1
X_542_ i_reg2_data[31] imm_i\[31\] op2_sel VSS VSS VCC VCC _166_ sky130_fd_sc_hd__mux2_1
X_809_ _354_ _359_ VSS VSS VCC VCC _360_ sky130_fd_sc_hd__and2_1
X_456_ _121_ VSS VSS VCC VCC o_op1[21] sky130_fd_sc_hd__buf_2
X_525_ _157_ VSS VSS VCC VCC o_op2[22] sky130_fd_sc_hd__buf_2
X_439_ i_reg1_data[13] o_pc[13] op1_sel VSS VSS VCC VCC _113_ sky130_fd_sc_hd__mux2_1
X_508_ _148_ VSS VSS VCC VCC o_op2[14] sky130_fd_sc_hd__buf_2
X_790_ i_inst_branch o_inst_branch _290_ VSS VSS VCC VCC _347_ sky130_fd_sc_hd__mux2_1
X_988_ clknet_3_6__leaf_i_clk _047_ VSS VSS VCC VCC o_pc_next[7] sky130_fd_sc_hd__dfxtp_2
X_842_ i_pc[4] o_pc[4] _379_ VSS VSS VCC VCC _380_ sky130_fd_sc_hd__mux2_1
X_911_ clknet_3_2__leaf_i_clk _067_ VSS VSS VCC VCC o_rs2[1] sky130_fd_sc_hd__dfxtp_2
X_773_ i_imm_i[28] imm_i\[28\] _328_ VSS VSS VCC VCC _337_ sky130_fd_sc_hd__mux2_1
X_825_ _370_ VSS VSS VCC VCC _020_ sky130_fd_sc_hd__clkbuf_1
X_756_ _280_ VSS VSS VCC VCC _328_ sky130_fd_sc_hd__clkbuf_4
X_687_ _288_ VSS VSS VCC VCC _289_ sky130_fd_sc_hd__buf_2
X_610_ _174_ VSS VSS VCC VCC _225_ sky130_fd_sc_hd__buf_2
X_472_ _129_ VSS VSS VCC VCC o_op1[29] sky130_fd_sc_hd__buf_2
X_541_ _165_ VSS VSS VCC VCC o_op2[30] sky130_fd_sc_hd__buf_2
X_808_ i_alu_ctrl[3] o_alu_ctrl[3] _351_ VSS VSS VCC VCC _359_ sky130_fd_sc_hd__mux2_1
X_739_ _319_ VSS VSS VCC VCC _082_ sky130_fd_sc_hd__clkbuf_1
X_455_ _097_ i_reg1_data[21] VSS VSS VCC VCC _121_ sky130_fd_sc_hd__and2b_1
X_524_ i_reg2_data[22] imm_i\[22\] _153_ VSS VSS VCC VCC _157_ sky130_fd_sc_hd__mux2_1
X_438_ _112_ VSS VSS VCC VCC o_op1[12] sky130_fd_sc_hd__buf_2
X_507_ i_reg2_data[14] imm_i\[14\] _142_ VSS VSS VCC VCC _148_ sky130_fd_sc_hd__mux2_1
X_987_ clknet_3_6__leaf_i_clk _046_ VSS VSS VCC VCC o_pc_next[6] sky130_fd_sc_hd__dfxtp_2
X_910_ clknet_3_2__leaf_i_clk _066_ VSS VSS VCC VCC o_rs2[0] sky130_fd_sc_hd__dfxtp_2
X_841_ _280_ VSS VSS VCC VCC _379_ sky130_fd_sc_hd__clkbuf_4
X_772_ _336_ VSS VSS VCC VCC _001_ sky130_fd_sc_hd__clkbuf_1
X_824_ _354_ _369_ VSS VSS VCC VCC _370_ sky130_fd_sc_hd__and2_1
X_755_ _327_ VSS VSS VCC VCC _090_ sky130_fd_sc_hd__clkbuf_1
X_686_ i_flush i_reset_n VSS VSS VCC VCC _288_ sky130_fd_sc_hd__and2b_1
X_540_ i_reg2_data[30] imm_i\[30\] op2_sel VSS VSS VCC VCC _165_ sky130_fd_sc_hd__mux2_1
X_471_ _099_ i_reg1_data[29] VSS VSS VCC VCC _129_ sky130_fd_sc_hd__and2b_1
X_807_ _358_ VSS VSS VCC VCC _014_ sky130_fd_sc_hd__clkbuf_1
X_669_ imm_i\[1\] i_ret_addr[1] _167_ VSS VSS VCC VCC _277_ sky130_fd_sc_hd__mux2_1
X_738_ i_imm_i[11] imm_i\[11\] _317_ VSS VSS VCC VCC _319_ sky130_fd_sc_hd__mux2_1
X_523_ _156_ VSS VSS VCC VCC o_op2[21] sky130_fd_sc_hd__buf_2
X_454_ _120_ VSS VSS VCC VCC o_op1[20] sky130_fd_sc_hd__buf_2
X_506_ _147_ VSS VSS VCC VCC o_op2[13] sky130_fd_sc_hd__buf_2
X_437_ i_reg1_data[12] o_pc[12] _102_ VSS VSS VCC VCC _112_ sky130_fd_sc_hd__mux2_1
X_986_ clknet_3_6__leaf_i_clk _045_ VSS VSS VCC VCC o_pc_next[5] sky130_fd_sc_hd__dfxtp_2
X_840_ _378_ VSS VSS VCC VCC _027_ sky130_fd_sc_hd__clkbuf_1
X_771_ i_imm_i[27] imm_i\[27\] _328_ VSS VSS VCC VCC _336_ sky130_fd_sc_hd__mux2_1
X_969_ clknet_3_0__leaf_i_clk _028_ VSS VSS VCC VCC o_pc[4] sky130_fd_sc_hd__dfxtp_4
X_823_ i_res_src[2] o_res_src[2] _351_ VSS VSS VCC VCC _369_ sky130_fd_sc_hd__mux2_1
X_754_ i_imm_i[19] imm_i\[19\] _317_ VSS VSS VCC VCC _327_ sky130_fd_sc_hd__mux2_1
X_685_ _287_ VSS VSS VCC VCC _060_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_3__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_3__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_470_ _128_ VSS VSS VCC VCC o_op1[28] sky130_fd_sc_hd__buf_2
X_806_ _354_ _357_ VSS VSS VCC VCC _358_ sky130_fd_sc_hd__and2_1
X_668_ _274_ _276_ VSS VSS VCC VCC o_pc_target[15] sky130_fd_sc_hd__xnor2_4
X_737_ _318_ VSS VSS VCC VCC _081_ sky130_fd_sc_hd__clkbuf_1
X_599_ _212_ _215_ VSS VSS VCC VCC o_pc_target[7] sky130_fd_sc_hd__xnor2_4
X_453_ _097_ i_reg1_data[20] VSS VSS VCC VCC _120_ sky130_fd_sc_hd__and2b_1
X_522_ i_reg2_data[21] imm_i\[21\] _153_ VSS VSS VCC VCC _156_ sky130_fd_sc_hd__mux2_1
X_436_ _111_ VSS VSS VCC VCC o_op1[11] sky130_fd_sc_hd__buf_2
X_505_ i_reg2_data[13] imm_i\[13\] _142_ VSS VSS VCC VCC _147_ sky130_fd_sc_hd__mux2_1
X_985_ clknet_3_3__leaf_i_clk _044_ VSS VSS VCC VCC o_pc_next[4] sky130_fd_sc_hd__dfxtp_2
X_419_ i_reg1_data[3] o_pc[3] _102_ VSS VSS VCC VCC _103_ sky130_fd_sc_hd__mux2_1
X_770_ _335_ VSS VSS VCC VCC _000_ sky130_fd_sc_hd__clkbuf_1
X_968_ clknet_3_0__leaf_i_clk _027_ VSS VSS VCC VCC o_pc[3] sky130_fd_sc_hd__dfxtp_2
X_899_ _409_ VSS VSS VCC VCC _055_ sky130_fd_sc_hd__clkbuf_1
X_822_ _368_ VSS VSS VCC VCC _019_ sky130_fd_sc_hd__clkbuf_1
X_753_ _326_ VSS VSS VCC VCC _089_ sky130_fd_sc_hd__clkbuf_1
X_684_ i_rs1[4] o_rs1[4] _282_ VSS VSS VCC VCC _287_ sky130_fd_sc_hd__mux2_1
X_805_ i_alu_ctrl[2] o_alu_ctrl[2] _351_ VSS VSS VCC VCC _357_ sky130_fd_sc_hd__mux2_1
X_736_ i_imm_i[10] imm_i\[10\] _317_ VSS VSS VCC VCC _318_ sky130_fd_sc_hd__mux2_1
X_667_ _266_ _275_ VSS VSS VCC VCC _276_ sky130_fd_sc_hd__or2_2
X_598_ _195_ _213_ _214_ VSS VSS VCC VCC _215_ sky130_fd_sc_hd__o21a_1
X_452_ _119_ VSS VSS VCC VCC o_op1[19] sky130_fd_sc_hd__buf_2
X_521_ _155_ VSS VSS VCC VCC o_op2[20] sky130_fd_sc_hd__buf_2
X_719_ i_imm_i[2] imm_i\[2\] _306_ VSS VSS VCC VCC _309_ sky130_fd_sc_hd__mux2_1
X_435_ i_reg1_data[11] o_pc[11] _102_ VSS VSS VCC VCC _111_ sky130_fd_sc_hd__mux2_1
X_504_ _146_ VSS VSS VCC VCC o_op2[12] sky130_fd_sc_hd__buf_2
X_984_ clknet_3_3__leaf_i_clk _043_ VSS VSS VCC VCC o_pc_next[3] sky130_fd_sc_hd__dfxtp_2
X_418_ op1_sel VSS VSS VCC VCC _102_ sky130_fd_sc_hd__clkbuf_4
X_898_ i_pc_next[15] o_pc_next[15] _281_ VSS VSS VCC VCC _409_ sky130_fd_sc_hd__mux2_1
X_967_ clknet_3_1__leaf_i_clk _026_ VSS VSS VCC VCC o_pc[2] sky130_fd_sc_hd__dfxtp_2
X_821_ _354_ _367_ VSS VSS VCC VCC _368_ sky130_fd_sc_hd__and2_1
X_752_ i_imm_i[18] imm_i\[18\] _317_ VSS VSS VCC VCC _326_ sky130_fd_sc_hd__mux2_1
X_683_ _286_ VSS VSS VCC VCC _059_ sky130_fd_sc_hd__clkbuf_1
X_804_ _356_ VSS VSS VCC VCC _013_ sky130_fd_sc_hd__clkbuf_1
X_735_ _281_ VSS VSS VCC VCC _317_ sky130_fd_sc_hd__clkbuf_4
X_666_ _259_ _263_ _267_ _269_ VSS VSS VCC VCC _275_ sky130_fd_sc_hd__a211oi_1
X_597_ imm_i\[6\] _203_ _205_ _197_ VSS VSS VCC VCC _214_ sky130_fd_sc_hd__a22oi_2
X_520_ i_reg2_data[20] imm_i\[20\] _153_ VSS VSS VCC VCC _155_ sky130_fd_sc_hd__mux2_1
X_451_ _097_ i_reg1_data[19] VSS VSS VCC VCC _119_ sky130_fd_sc_hd__and2b_1
X_649_ _245_ _253_ VSS VSS VCC VCC _260_ sky130_fd_sc_hd__nand2_1
X_718_ _308_ VSS VSS VCC VCC _072_ sky130_fd_sc_hd__clkbuf_1
X_503_ i_reg2_data[12] imm_i\[12\] _142_ VSS VSS VCC VCC _146_ sky130_fd_sc_hd__mux2_1
X_434_ _110_ VSS VSS VCC VCC o_op1[10] sky130_fd_sc_hd__buf_2
X_983_ clknet_3_3__leaf_i_clk _042_ VSS VSS VCC VCC o_pc_next[2] sky130_fd_sc_hd__dfxtp_2
X_417_ _101_ VSS VSS VCC VCC o_op1[2] sky130_fd_sc_hd__buf_2
X_897_ _408_ VSS VSS VCC VCC _054_ sky130_fd_sc_hd__clkbuf_1
X_966_ clknet_3_1__leaf_i_clk _025_ VSS VSS VCC VCC o_pc[1] sky130_fd_sc_hd__dfxtp_2
X_820_ i_res_src[1] o_res_src[1] _351_ VSS VSS VCC VCC _367_ sky130_fd_sc_hd__mux2_1
X_751_ _325_ VSS VSS VCC VCC _088_ sky130_fd_sc_hd__clkbuf_1
X_682_ i_rs1[3] o_rs1[3] _282_ VSS VSS VCC VCC _286_ sky130_fd_sc_hd__mux2_1
X_949_ clknet_3_5__leaf_i_clk _008_ VSS VSS VCC VCC inst_jal sky130_fd_sc_hd__dfxtp_1
X_803_ _354_ _355_ VSS VSS VCC VCC _356_ sky130_fd_sc_hd__and2_1
X_665_ _167_ i_ret_addr[15] _272_ _273_ VSS VSS VCC VCC _274_ sky130_fd_sc_hd__a22o_2
X_734_ _316_ VSS VSS VCC VCC _080_ sky130_fd_sc_hd__clkbuf_1
X_596_ _200_ _206_ VSS VSS VCC VCC _213_ sky130_fd_sc_hd__nand2_1
X_450_ _118_ VSS VSS VCC VCC o_op1[18] sky130_fd_sc_hd__buf_2
X_648_ _255_ _256_ _258_ VSS VSS VCC VCC _259_ sky130_fd_sc_hd__mux2_2
X_717_ i_imm_i[1] imm_i\[1\] _306_ VSS VSS VCC VCC _308_ sky130_fd_sc_hd__mux2_1
X_579_ imm_i\[5\] i_ret_addr[5] inst_mret VSS VSS VCC VCC _198_ sky130_fd_sc_hd__mux2_1
X_433_ i_reg1_data[10] o_pc[10] _102_ VSS VSS VCC VCC _110_ sky130_fd_sc_hd__mux2_1
X_502_ _145_ VSS VSS VCC VCC o_op2[11] sky130_fd_sc_hd__buf_2
X_982_ clknet_3_3__leaf_i_clk _041_ VSS VSS VCC VCC o_pc_next[1] sky130_fd_sc_hd__dfxtp_2
X_416_ i_reg1_data[2] o_pc[2] _099_ VSS VSS VCC VCC _101_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_6__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_965_ clknet_3_5__leaf_i_clk _024_ VSS VSS VCC VCC o_funct3[2] sky130_fd_sc_hd__dfxtp_2
X_896_ i_pc_next[14] o_pc_next[14] _281_ VSS VSS VCC VCC _408_ sky130_fd_sc_hd__mux2_1
X_750_ i_imm_i[17] imm_i\[17\] _317_ VSS VSS VCC VCC _325_ sky130_fd_sc_hd__mux2_1
X_681_ _285_ VSS VSS VCC VCC _058_ sky130_fd_sc_hd__clkbuf_1
X_948_ clknet_3_5__leaf_i_clk _007_ VSS VSS VCC VCC inst_jalr sky130_fd_sc_hd__dfxtp_4
X_879_ _399_ VSS VSS VCC VCC _045_ sky130_fd_sc_hd__clkbuf_1
X_802_ i_alu_ctrl[1] o_alu_ctrl[1] _351_ VSS VSS VCC VCC _355_ sky130_fd_sc_hd__mux2_1
X_664_ imm_i\[15\] _271_ _167_ VSS VSS VCC VCC _273_ sky130_fd_sc_hd__a21oi_1
X_733_ i_imm_i[9] imm_i\[9\] _306_ VSS VSS VCC VCC _316_ sky130_fd_sc_hd__mux2_1
X_595_ _209_ _211_ VSS VSS VCC VCC _212_ sky130_fd_sc_hd__nor2_2
X_716_ _307_ VSS VSS VCC VCC _071_ sky130_fd_sc_hd__clkbuf_1
X_647_ _225_ _257_ VSS VSS VCC VCC _258_ sky130_fd_sc_hd__nand2_1
X_578_ _174_ imm_i\[5\] _196_ VSS VSS VCC VCC _197_ sky130_fd_sc_hd__and3_1
