
.include ../block_head.spice
.include simulation/pc_inc.spice

.include simulation/stimuli_pc_inc.cir

.tran 100p 14n
.print tran format=raw file=simulation/pc_inc.spice.raw v(*)

.end
