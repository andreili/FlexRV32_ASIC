magic
tech sky130A
magscale 1 2
timestamp 1684682343
<< nwell >>
rect 80 230 1875 505
<< pwell >>
rect 80 -130 1875 45
<< nmos >>
rect 185 -90 215 5
rect 280 -90 310 5
rect 495 -90 525 5
rect 630 -90 660 5
rect 775 -90 805 5
rect 910 -90 940 5
rect 1005 -90 1035 5
rect 1150 -90 1180 5
rect 1295 -90 1325 5
rect 1430 -90 1460 5
rect 1525 -90 1555 5
rect 1740 -90 1770 5
<< pmos >>
rect 185 270 215 465
rect 280 270 310 465
rect 495 270 525 465
rect 630 270 660 465
rect 775 270 805 465
rect 910 270 940 465
rect 1005 270 1035 465
rect 1150 270 1180 465
rect 1295 270 1325 465
rect 1430 270 1460 465
rect 1525 270 1555 465
rect 1740 270 1770 465
<< ndiff >>
rect 120 -5 185 5
rect 120 -40 135 -5
rect 170 -40 185 -5
rect 120 -90 185 -40
rect 215 -45 280 5
rect 215 -80 230 -45
rect 265 -80 280 -45
rect 215 -90 280 -80
rect 310 -5 375 5
rect 310 -40 325 -5
rect 360 -40 375 -5
rect 310 -90 375 -40
rect 430 -45 495 5
rect 430 -80 445 -45
rect 480 -80 495 -45
rect 430 -90 495 -80
rect 525 -5 630 5
rect 525 -40 560 -5
rect 595 -40 630 -5
rect 525 -90 630 -40
rect 660 -5 775 5
rect 660 -40 700 -5
rect 735 -40 775 -5
rect 660 -90 775 -40
rect 805 -5 910 5
rect 805 -40 840 -5
rect 875 -40 910 -5
rect 805 -90 910 -40
rect 940 -45 1005 5
rect 940 -80 955 -45
rect 990 -80 1005 -45
rect 940 -90 1005 -80
rect 1035 -5 1150 5
rect 1035 -40 1075 -5
rect 1110 -40 1150 -5
rect 1035 -90 1150 -40
rect 1180 -5 1295 5
rect 1180 -40 1220 -5
rect 1255 -40 1295 -5
rect 1180 -90 1295 -40
rect 1325 -5 1430 5
rect 1325 -40 1360 -5
rect 1395 -40 1430 -5
rect 1325 -90 1430 -40
rect 1460 -45 1525 5
rect 1460 -80 1475 -45
rect 1510 -80 1525 -45
rect 1460 -90 1525 -80
rect 1555 -5 1620 5
rect 1555 -40 1570 -5
rect 1605 -40 1620 -5
rect 1555 -90 1620 -40
rect 1675 -45 1740 5
rect 1675 -80 1690 -45
rect 1725 -80 1740 -45
rect 1675 -90 1740 -80
rect 1770 -5 1835 5
rect 1770 -40 1785 -5
rect 1820 -40 1835 -5
rect 1770 -90 1835 -40
<< pdiff >>
rect 120 315 185 465
rect 120 280 135 315
rect 170 280 185 315
rect 120 270 185 280
rect 215 455 280 465
rect 215 420 230 455
rect 265 420 280 455
rect 215 270 280 420
rect 310 315 375 465
rect 310 280 325 315
rect 360 280 375 315
rect 310 270 375 280
rect 430 455 495 465
rect 430 420 445 455
rect 480 420 495 455
rect 430 270 495 420
rect 525 315 630 465
rect 525 280 560 315
rect 595 280 630 315
rect 525 270 630 280
rect 660 315 775 465
rect 660 280 700 315
rect 735 280 775 315
rect 660 270 775 280
rect 805 315 910 465
rect 805 280 840 315
rect 875 280 910 315
rect 805 270 910 280
rect 940 455 1005 465
rect 940 420 955 455
rect 990 420 1005 455
rect 940 270 1005 420
rect 1035 315 1150 465
rect 1035 280 1075 315
rect 1110 280 1150 315
rect 1035 270 1150 280
rect 1180 315 1295 465
rect 1180 280 1220 315
rect 1255 280 1295 315
rect 1180 270 1295 280
rect 1325 315 1430 465
rect 1325 280 1360 315
rect 1395 280 1430 315
rect 1325 270 1430 280
rect 1460 455 1525 465
rect 1460 420 1475 455
rect 1510 420 1525 455
rect 1460 270 1525 420
rect 1555 315 1620 465
rect 1555 280 1570 315
rect 1605 280 1620 315
rect 1555 270 1620 280
rect 1675 455 1740 465
rect 1675 420 1690 455
rect 1725 420 1740 455
rect 1675 270 1740 420
rect 1770 315 1835 465
rect 1770 280 1785 315
rect 1820 280 1835 315
rect 1770 270 1835 280
<< ndiffc >>
rect 135 -40 170 -5
rect 230 -80 265 -45
rect 325 -40 360 -5
rect 445 -80 480 -45
rect 560 -40 595 -5
rect 700 -40 735 -5
rect 840 -40 875 -5
rect 955 -80 990 -45
rect 1075 -40 1110 -5
rect 1220 -40 1255 -5
rect 1360 -40 1395 -5
rect 1475 -80 1510 -45
rect 1570 -40 1605 -5
rect 1690 -80 1725 -45
rect 1785 -40 1820 -5
<< pdiffc >>
rect 135 280 170 315
rect 230 420 265 455
rect 325 280 360 315
rect 445 420 480 455
rect 560 280 595 315
rect 700 280 735 315
rect 840 280 875 315
rect 955 420 990 455
rect 1075 280 1110 315
rect 1220 280 1255 315
rect 1360 280 1395 315
rect 1475 420 1510 455
rect 1570 280 1605 315
rect 1690 420 1725 455
rect 1785 280 1820 315
<< poly >>
rect 185 465 215 495
rect 280 465 310 495
rect 495 465 525 495
rect 630 465 660 495
rect 775 465 805 495
rect 910 465 940 495
rect 1005 465 1035 495
rect 1150 465 1180 495
rect 1295 465 1325 495
rect 1430 465 1460 495
rect 1525 465 1555 495
rect 1740 465 1770 495
rect 185 235 215 270
rect 180 215 235 235
rect 180 180 190 215
rect 225 180 235 215
rect 180 160 235 180
rect 185 5 215 160
rect 280 115 310 270
rect 495 235 525 270
rect 630 235 660 270
rect 775 235 805 270
rect 405 215 525 235
rect 405 180 415 215
rect 450 180 525 215
rect 405 160 525 180
rect 620 215 675 235
rect 620 180 630 215
rect 665 180 675 215
rect 620 160 675 180
rect 760 215 815 235
rect 760 180 770 215
rect 805 180 815 215
rect 760 160 815 180
rect 260 95 315 115
rect 260 60 270 95
rect 305 60 315 95
rect 260 40 315 60
rect 280 5 310 40
rect 495 5 525 160
rect 910 115 940 270
rect 1005 235 1035 270
rect 1150 235 1180 270
rect 1295 235 1325 270
rect 995 215 1050 235
rect 995 180 1005 215
rect 1040 180 1050 215
rect 995 160 1050 180
rect 1140 215 1195 235
rect 1140 180 1150 215
rect 1185 180 1195 215
rect 1140 160 1195 180
rect 1280 215 1335 235
rect 1280 180 1290 215
rect 1325 180 1335 215
rect 1430 205 1460 270
rect 1280 160 1335 180
rect 1420 185 1475 205
rect 585 105 660 115
rect 585 70 605 105
rect 640 70 660 105
rect 585 60 660 70
rect 630 5 660 60
rect 760 95 815 115
rect 760 60 770 95
rect 805 60 815 95
rect 760 40 815 60
rect 900 95 955 115
rect 900 60 910 95
rect 945 60 955 95
rect 900 40 955 60
rect 775 5 805 40
rect 910 5 940 40
rect 1005 5 1035 160
rect 1420 150 1430 185
rect 1465 150 1475 185
rect 1420 130 1475 150
rect 1140 95 1195 115
rect 1140 60 1150 95
rect 1185 60 1195 95
rect 1140 40 1195 60
rect 1280 95 1335 115
rect 1280 60 1290 95
rect 1325 60 1335 95
rect 1280 40 1335 60
rect 1150 5 1180 40
rect 1295 5 1325 40
rect 1430 5 1460 130
rect 1525 115 1555 270
rect 1525 95 1580 115
rect 1740 110 1770 270
rect 1525 60 1535 95
rect 1570 60 1580 95
rect 1525 40 1580 60
rect 1695 90 1770 110
rect 1695 55 1705 90
rect 1740 55 1770 90
rect 1525 5 1555 40
rect 1695 35 1770 55
rect 1740 5 1770 35
rect 185 -120 215 -90
rect 280 -120 310 -90
rect 495 -120 525 -90
rect 630 -120 660 -90
rect 775 -120 805 -90
rect 910 -120 940 -90
rect 1005 -120 1035 -90
rect 1150 -120 1180 -90
rect 1295 -120 1325 -90
rect 1430 -120 1460 -90
rect 1525 -120 1555 -90
rect 1740 -120 1770 -90
<< polycont >>
rect 190 180 225 215
rect 415 180 450 215
rect 630 180 665 215
rect 770 180 805 215
rect 270 60 305 95
rect 1005 180 1040 215
rect 1150 180 1185 215
rect 1290 180 1325 215
rect 605 70 640 105
rect 770 60 805 95
rect 910 60 945 95
rect 1430 150 1465 185
rect 1150 60 1185 95
rect 1290 60 1325 95
rect 1535 60 1570 95
rect 1705 55 1740 90
<< locali >>
rect 120 470 1835 520
rect 230 455 265 470
rect 230 400 265 420
rect 445 455 480 470
rect 445 400 480 420
rect 955 455 990 470
rect 955 400 990 420
rect 1475 455 1510 470
rect 1475 400 1510 420
rect 1690 455 1725 470
rect 1690 400 1725 420
rect 120 315 190 335
rect 120 280 135 315
rect 170 280 190 315
rect 120 270 190 280
rect 305 315 380 335
rect 305 280 325 315
rect 360 280 380 315
rect 305 270 380 280
rect 120 115 155 270
rect 190 215 235 235
rect 225 180 235 215
rect 190 160 235 180
rect 120 95 305 115
rect 120 60 270 95
rect 120 40 305 60
rect 120 5 155 40
rect 120 -5 190 5
rect 340 -5 380 270
rect 495 315 595 335
rect 495 280 560 315
rect 495 245 595 280
rect 700 315 735 335
rect 415 215 460 235
rect 450 180 460 215
rect 415 160 460 180
rect 495 30 530 245
rect 630 215 665 235
rect 630 160 665 180
rect 585 105 660 115
rect 585 70 605 105
rect 640 70 660 105
rect 585 65 660 70
rect 495 -5 595 30
rect 120 -40 135 -5
rect 170 -40 190 -5
rect 120 -60 190 -40
rect 230 -45 265 -25
rect 305 -40 325 -5
rect 360 -40 380 -5
rect 540 -40 560 -5
rect 230 -95 265 -80
rect 425 -80 445 -45
rect 480 -80 500 -45
rect 540 -60 595 -40
rect 700 -5 735 280
rect 840 315 875 335
rect 770 215 805 235
rect 770 160 805 180
rect 700 -60 735 -40
rect 770 95 805 115
rect 770 -5 805 60
rect 770 -60 805 -40
rect 840 -5 875 280
rect 940 315 1040 335
rect 940 280 950 315
rect 985 280 1040 315
rect 940 215 1040 280
rect 940 180 1005 215
rect 940 160 1040 180
rect 1075 315 1110 335
rect 1075 115 1110 280
rect 1150 315 1185 335
rect 1150 215 1185 280
rect 1150 160 1185 180
rect 1220 315 1255 335
rect 1785 315 1820 335
rect 910 95 1110 115
rect 945 60 1110 95
rect 910 40 1110 60
rect 1075 -5 1110 40
rect 840 -60 875 -40
rect 955 -45 990 -25
rect 425 -95 500 -80
rect 1075 -60 1110 -40
rect 1150 95 1185 115
rect 1150 -5 1185 60
rect 1150 -60 1185 -40
rect 1220 5 1255 280
rect 1340 280 1360 315
rect 1395 280 1415 315
rect 1340 270 1415 280
rect 1550 280 1570 315
rect 1605 280 1645 315
rect 1550 275 1645 280
rect 1290 215 1325 235
rect 1290 160 1325 180
rect 1290 95 1325 115
rect 1290 40 1325 60
rect 1360 5 1395 270
rect 1430 185 1475 205
rect 1605 185 1645 275
rect 1465 150 1645 185
rect 1430 130 1475 150
rect 1520 95 1570 115
rect 1520 60 1535 95
rect 1520 40 1570 60
rect 1605 110 1645 150
rect 1605 90 1745 110
rect 1605 55 1705 90
rect 1740 55 1745 90
rect 1605 35 1745 55
rect 1220 -5 1305 5
rect 1290 -40 1305 -5
rect 1340 -5 1415 5
rect 1605 0 1645 35
rect 1340 -40 1360 -5
rect 1395 -40 1415 -5
rect 1550 -5 1645 0
rect 1220 -60 1305 -40
rect 1475 -45 1510 -25
rect 1550 -40 1570 -5
rect 1605 -40 1645 -5
rect 1785 -5 1820 280
rect 955 -95 990 -80
rect 1475 -95 1510 -80
rect 1690 -45 1725 -25
rect 1785 -60 1820 -40
rect 1690 -95 1725 -80
rect 120 -145 1835 -95
<< viali >>
rect 270 60 305 95
rect 700 280 735 315
rect 630 180 665 215
rect 605 70 640 105
rect 325 -40 360 -5
rect 770 180 805 215
rect 770 -40 805 -5
rect 950 280 985 315
rect 1150 280 1185 315
rect 1150 -40 1185 -5
rect 1290 180 1325 215
rect 1290 60 1325 95
rect 1535 60 1570 95
rect 1255 -40 1290 -5
<< metal1 >>
rect 495 355 1105 410
rect 495 115 560 355
rect 1040 325 1105 355
rect 685 315 1000 325
rect 685 280 700 315
rect 735 280 950 315
rect 985 280 1000 315
rect 685 270 1000 280
rect 1040 315 1435 325
rect 1040 280 1150 315
rect 1185 280 1435 315
rect 1040 270 1435 280
rect 1040 235 1105 270
rect 1005 230 1105 235
rect 615 215 730 225
rect 615 180 630 215
rect 665 180 730 215
rect 615 170 730 180
rect 690 125 730 170
rect 760 215 1105 230
rect 760 180 770 215
rect 805 180 1105 215
rect 760 160 1105 180
rect 1135 215 1340 225
rect 1135 180 1290 215
rect 1325 180 1340 215
rect 1135 170 1340 180
rect 255 105 655 115
rect 255 95 605 105
rect 255 60 270 95
rect 305 70 605 95
rect 640 70 655 105
rect 305 60 655 70
rect 690 60 805 125
rect 255 50 655 60
rect 750 5 805 60
rect 1135 5 1200 170
rect 1380 105 1435 270
rect 1275 95 1435 105
rect 1275 60 1290 95
rect 1325 60 1435 95
rect 1275 50 1435 60
rect 1520 95 1580 115
rect 1520 60 1535 95
rect 1570 60 1580 95
rect 1520 5 1580 60
rect 305 -5 1200 5
rect 305 -40 325 -5
rect 360 -40 770 -5
rect 805 -40 1150 -5
rect 1185 -40 1200 -5
rect 305 -50 1200 -40
rect 1240 -5 1580 5
rect 1240 -40 1255 -5
rect 1290 -40 1580 -5
rect 1240 -50 1580 -40
<< labels >>
flabel locali 415 180 450 215 5 FreeSans 200 0 0 0 i_data
port 1 nsew signal input
flabel locali 190 180 225 215 5 FreeSans 200 0 0 0 i_clk
port 2 nsew signal input
flabel locali 1785 55 1820 90 5 FreeSans 200 0 0 0 Qp
port 3 nsew signal output
flabel locali 1705 55 1740 90 5 FreeSans 200 0 0 0 Qn
port 4 nsew signal output
flabel locali 135 -135 170 -100 5 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali 135 475 170 510 5 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel pwell 135 -135 170 -100 5 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell 135 475 170 510 5 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel locali 120 5 155 30 5 pcb
rlabel locali 340 5 375 30 5 pc
rlabel locali 560 5 595 30 5 db
rlabel locali 700 5 735 30 5 db1
rlabel locali 840 5 875 30 5 db1l
rlabel locali 1075 5 1110 30 5 db1b
rlabel locali 1220 5 1255 30 5 db2
rlabel locali 1360 5 1395 30 5 db2l
<< end >>
