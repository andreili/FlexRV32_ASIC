* NGSPICE file created from rv_decode.ext - technology: sky130A


X_0985_ clknet_3_1_0_i_clk _0026_ VSS VSS VCC VCC o_rd[3] sky130_fd_sc_hd__dfxtp_2
X_0770_ _0170_ _0198_ _0163_ i_instruction[12] VSS VSS VCC VCC _0297_ sky130_fd_sc_hd__and4b_2
X_0968_ clknet_3_7_0_i_clk _0009_ VSS VSS VCC VCC o_csr_pc_next[10] sky130_fd_sc_hd__dfxtp_2
X_0899_ _0166_ _0240_ _0242_ _0329_ i_instruction[3] VSS VSS VCC VCC _0411_
+ sky130_fd_sc_hd__a32o_1
X_0822_ _0272_ _0285_ _0297_ _0337_ VSS VSS VCC VCC _0343_ sky130_fd_sc_hd__a211o_1
X_0753_ i_instruction[4] _0250_ _0274_ i_instruction[9] _0248_ VSS VSS VCC VCC
+ _0283_ sky130_fd_sc_hd__a221o_1
X_0684_ _0164_ _0170_ VSS VSS VCC VCC _0219_ sky130_fd_sc_hd__nand2_4
X_1021_ clknet_3_1_0_i_clk _0062_ VSS VSS VCC VCC o_pc[15] sky130_fd_sc_hd__dfxtp_2
X_0805_ _0172_ _0327_ _0208_ VSS VSS VCC VCC _0328_ sky130_fd_sc_hd__o21a_1
X_0736_ _0183_ VSS VSS VCC VCC _0267_ sky130_fd_sc_hd__inv_2
X_0667_ _0196_ _0203_ i_stall VSS VSS VCC VCC _0204_ sky130_fd_sc_hd__a21o_1
X_0598_ o_csr_pc_next[7] i_pc_next[7] _0140_ VSS VSS VCC VCC _0147_ sky130_fd_sc_hd__mux2_1
X_0521_ _0111_ VSS VSS VCC VCC o_imm_i[6] sky130_fd_sc_hd__buf_2
X_0452_ instruction\[4\] VSS VSS VCC VCC _0064_ sky130_fd_sc_hd__clkinv_2
X_1004_ clknet_3_6_0_i_clk _0045_ VSS VSS VCC VCC o_csr_idx[9] sky130_fd_sc_hd__dfxtp_4
X_0719_ _0246_ _0219_ _0189_ VSS VSS VCC VCC _0251_ sky130_fd_sc_hd__o21a_1
X_0504_ _0100_ VSS VSS VCC VCC _0101_ sky130_fd_sc_hd__buf_12
X_0984_ clknet_3_4_0_i_clk _0025_ VSS VSS VCC VCC o_rd[2] sky130_fd_sc_hd__dfxtp_2
X_0967_ clknet_3_7_0_i_clk _0008_ VSS VSS VCC VCC o_csr_pc_next[9] sky130_fd_sc_hd__dfxtp_2
X_0898_ _0349_ o_csr_idx[6] _0313_ _0410_ VSS VSS VCC VCC _0042_ sky130_fd_sc_hd__o211a_1
X_0821_ _0158_ o_csr_imm[2] _0340_ _0342_ _0216_ VSS VSS VCC VCC _0033_ sky130_fd_sc_hd__o221a_1
X_0752_ _0281_ _0270_ _0195_ VSS VSS VCC VCC _0282_ sky130_fd_sc_hd__o21a_1
X_0683_ i_instruction[4] _0206_ _0184_ VSS VSS VCC VCC _0218_ sky130_fd_sc_hd__a21o_1
X_1020_ clknet_3_2_0_i_clk _0061_ VSS VSS VCC VCC o_pc[14] sky130_fd_sc_hd__dfxtp_2
X_0804_ _0189_ _0318_ _0177_ VSS VSS VCC VCC _0327_ sky130_fd_sc_hd__o21a_1
X_0735_ i_instruction[1] _0177_ _0265_ _0162_ VSS VSS VCC VCC _0266_ sky130_fd_sc_hd__a31o_1
X_0666_ _0202_ VSS VSS VCC VCC _0203_ sky130_fd_sc_hd__buf_4
X_0597_ _0146_ VSS VSS VCC VCC _0005_ sky130_fd_sc_hd__clkbuf_1
X_0520_ o_csr_idx[6] _0086_ VSS VSS VCC VCC _0111_ sky130_fd_sc_hd__and2_1
X_0451_ instruction\[3\] instruction\[2\] VSS VSS VCC VCC _0063_ sky130_fd_sc_hd__nor2_2
X_1003_ clknet_3_6_0_i_clk _0044_ VSS VSS VCC VCC o_csr_idx[8] sky130_fd_sc_hd__dfxtp_4
X_0718_ _0222_ VSS VSS VCC VCC _0250_ sky130_fd_sc_hd__buf_4
X_0649_ _0185_ _0186_ i_flush VSS VSS VCC VCC _0017_ sky130_fd_sc_hd__a21oi_1
X_0503_ _0068_ _0099_ VSS VSS VCC VCC _0100_ sky130_fd_sc_hd__or2_1
X_0983_ clknet_3_2_0_i_clk _0024_ VSS VSS VCC VCC o_rd[1] sky130_fd_sc_hd__dfxtp_2
X_0966_ clknet_3_0_0_i_clk _0007_ VSS VSS VCC VCC o_csr_pc_next[8] sky130_fd_sc_hd__dfxtp_2
X_0897_ _0162_ _0409_ VSS VSS VCC VCC _0410_ sky130_fd_sc_hd__or2_1
X_0820_ _0227_ _0341_ _0238_ VSS VSS VCC VCC _0342_ sky130_fd_sc_hd__a21o_1
X_0751_ _0165_ i_instruction[9] VSS VSS VCC VCC _0281_ sky130_fd_sc_hd__and2_1
X_0682_ _0159_ instruction\[3\] _0161_ _0217_ VSS VSS VCC VCC _0019_ sky130_fd_sc_hd__o211a_1
X_0949_ o_pc[11] i_pc[11] _0440_ VSS VSS VCC VCC _0446_ sky130_fd_sc_hd__mux2_1
X_0803_ _0159_ o_csr_imm[0] _0313_ _0326_ VSS VSS VCC VCC _0031_ sky130_fd_sc_hd__o211a_1
X_0734_ _0219_ _0213_ _0189_ i_instruction[0] VSS VSS VCC VCC _0265_ sky130_fd_sc_hd__a211o_1
X_0665_ _0170_ _0198_ i_ready VSS VSS VCC VCC _0202_ sky130_fd_sc_hd__and3b_1
X_0596_ o_csr_pc_next[6] i_pc_next[6] _0140_ VSS VSS VCC VCC _0146_ sky130_fd_sc_hd__mux2_1
X_1002_ clknet_3_2_0_i_clk _0043_ VSS VSS VCC VCC o_csr_idx[7] sky130_fd_sc_hd__dfxtp_2
X_0717_ _0247_ _0248_ _0195_ VSS VSS VCC VCC _0249_ sky130_fd_sc_hd__a21boi_1
X_0648_ _0168_ instruction\[1\] VSS VSS VCC VCC _0186_ sky130_fd_sc_hd__nand2_1
X_0579_ _0074_ _0134_ o_csr_read VSS VSS VCC VCC _0135_ sky130_fd_sc_hd__o21bai_4
X_0502_ _0098_ VSS VSS VCC VCC _0099_ sky130_fd_sc_hd__buf_2
X_0982_ clknet_3_4_0_i_clk _0023_ VSS VSS VCC VCC o_rd[0] sky130_fd_sc_hd__dfxtp_4
X_0965_ clknet_3_1_0_i_clk _0006_ VSS VSS VCC VCC o_csr_pc_next[7] sky130_fd_sc_hd__dfxtp_2
X_0896_ _0405_ _0407_ _0408_ _0244_ VSS VSS VCC VCC _0409_ sky130_fd_sc_hd__o22a_1
X_0750_ _0241_ _0213_ _0174_ VSS VSS VCC VCC _0280_ sky130_fd_sc_hd__o21ba_2
X_0681_ i_instruction[3] _0194_ _0204_ VSS VSS VCC VCC _0217_ sky130_fd_sc_hd__a21o_1
X_0948_ _0445_ VSS VSS VCC VCC _0057_ sky130_fd_sc_hd__clkbuf_1
X_0879_ _0242_ _0329_ i_instruction[2] VSS VSS VCC VCC _0393_ sky130_fd_sc_hd__o21a_1
X_0802_ _0181_ _0230_ _0320_ _0325_ VSS VSS VCC VCC _0326_ sky130_fd_sc_hd__a211o_1
X_0733_ _0158_ o_rd[0] _0260_ _0264_ _0216_ VSS VSS VCC VCC _0023_ sky130_fd_sc_hd__o221a_1
X_0664_ _0200_ VSS VSS VCC VCC _0201_ sky130_fd_sc_hd__inv_2
X_0595_ _0145_ VSS VSS VCC VCC _0004_ sky130_fd_sc_hd__clkbuf_1
X_1001_ clknet_3_6_0_i_clk _0042_ VSS VSS VCC VCC o_csr_idx[6] sky130_fd_sc_hd__dfxtp_4
X_0716_ _0170_ i_instruction[15] _0198_ _0163_ VSS VSS VCC VCC _0248_ sky130_fd_sc_hd__o31ai_4
X_0647_ _0169_ _0185_ i_flush VSS VSS VCC VCC _0016_ sky130_fd_sc_hd__a21oi_1
X_0578_ instruction\[4\] _0076_ _0085_ _0132_ _0133_ VSS VSS VCC VCC _0134_
+ sky130_fd_sc_hd__o41a_1
X_0501_ instruction\[4\] _0076_ instruction\[2\] VSS VSS VCC VCC _0098_ sky130_fd_sc_hd__and3_1
X_0981_ clknet_3_0_0_i_clk _0022_ VSS VSS VCC VCC instruction\[6\] sky130_fd_sc_hd__dfxtp_4
X_0964_ clknet_3_0_0_i_clk _0005_ VSS VSS VCC VCC o_csr_pc_next[6] sky130_fd_sc_hd__dfxtp_2
X_0895_ i_instruction[5] _0219_ _0256_ i_instruction[26] _0258_ vssd1 vssd1 vccd1
+ vccd1 _0408_ sky130_fd_sc_hd__o221a_1
Xclkbuf_3_6_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_6_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0680_ _0158_ instruction\[2\] _0205_ _0215_ _0216_ VSS VSS VCC VCC _0018_
+ sky130_fd_sc_hd__o221a_1
X_0947_ o_pc[10] i_pc[10] _0440_ VSS VSS VCC VCC _0445_ sky130_fd_sc_hd__mux2_1
X_0878_ _0158_ o_csr_idx[4] _0389_ _0392_ _0161_ VSS VSS VCC VCC _0040_ sky130_fd_sc_hd__o221a_1
X_0801_ _0249_ _0323_ _0324_ i_stall VSS VSS VCC VCC _0325_ sky130_fd_sc_hd__a211o_1
X_0732_ _0227_ _0263_ _0238_ VSS VSS VCC VCC _0264_ sky130_fd_sc_hd__a21o_1
X_0663_ _0197_ _0178_ _0199_ VSS VSS VCC VCC _0200_ sky130_fd_sc_hd__o21ai_4
X_0594_ o_csr_pc_next[5] i_pc_next[5] _0140_ VSS VSS VCC VCC _0145_ sky130_fd_sc_hd__mux2_1
X_1000_ clknet_3_3_0_i_clk _0041_ VSS VSS VCC VCC o_csr_idx[5] sky130_fd_sc_hd__dfxtp_4
X_0715_ _0165_ _0246_ VSS VSS VCC VCC _0247_ sky130_fd_sc_hd__nand2_1
X_0646_ _0172_ _0184_ _0158_ VSS VSS VCC VCC _0185_ sky130_fd_sc_hd__o21ai_1
X_0577_ _0064_ instruction\[2\] instruction\[3\] instruction\[6\] vssd1 vssd1 vccd1
+ vccd1 _0133_ sky130_fd_sc_hd__a211o_1
X_0500_ o_rd[0] o_inst_store _0096_ o_csr_idx[0] VSS VSS VCC VCC _0097_ sky130_fd_sc_hd__a22oi_2
X_0629_ _0162_ VSS VSS VCC VCC _0168_ sky130_fd_sc_hd__buf_6
Xclkbuf_0_i_clk i_clk VSS VSS VCC VCC clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_0980_ clknet_3_0_0_i_clk _0021_ VSS VSS VCC VCC instruction\[5\] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_3_2_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_2_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0963_ clknet_3_7_0_i_clk _0004_ VSS VSS VCC VCC o_csr_pc_next[5] sky130_fd_sc_hd__dfxtp_2
X_0894_ i_instruction[26] _0192_ _0207_ _0406_ _0187_ VSS VSS VCC VCC _0407_
+ sky130_fd_sc_hd__a221o_1
X_0946_ _0444_ VSS VSS VCC VCC _0056_ sky130_fd_sc_hd__clkbuf_1
X_0877_ _0166_ _0227_ _0390_ _0391_ VSS VSS VCC VCC _0392_ sky130_fd_sc_hd__a31o_1
X_0800_ _0246_ _0219_ _0311_ VSS VSS VCC VCC _0324_ sky130_fd_sc_hd__o21a_1
X_0731_ _0183_ _0210_ _0262_ VSS VSS VCC VCC _0263_ sky130_fd_sc_hd__a21o_1
X_0662_ i_instruction[15] _0198_ i_ready i_instruction[14] VSS VSS VCC VCC
+ _0199_ sky130_fd_sc_hd__and4b_2
X_0593_ _0144_ VSS VSS VCC VCC _0003_ sky130_fd_sc_hd__clkbuf_1
X_0929_ _0435_ VSS VSS VCC VCC _0048_ sky130_fd_sc_hd__clkbuf_1
X_0714_ i_instruction[7] VSS VSS VCC VCC _0246_ sky130_fd_sc_hd__buf_4
X_0645_ _0175_ _0183_ VSS VSS VCC VCC _0184_ sky130_fd_sc_hd__or2_1
X_0576_ o_csr_imm_sel o_funct3[1] instruction\[6\] instruction\[5\] vssd1 vssd1 vccd1
+ vccd1 _0132_ sky130_fd_sc_hd__or4_1
X_0628_ _0159_ valid_input _0161_ _0167_ VSS VSS VCC VCC _0015_ sky130_fd_sc_hd__o211a_1
X_0559_ o_csr_idx[5] _0072_ VSS VSS VCC VCC _0123_ sky130_fd_sc_hd__and2_1
X_0962_ clknet_3_4_0_i_clk _0003_ VSS VSS VCC VCC o_csr_pc_next[4] sky130_fd_sc_hd__dfxtp_2
X_0893_ i_instruction[2] _0261_ _0222_ _0246_ VSS VSS VCC VCC _0406_ sky130_fd_sc_hd__a22o_1
X_0945_ o_pc[9] i_pc[9] _0440_ VSS VSS VCC VCC _0444_ sky130_fd_sc_hd__mux2_1
X_0876_ i_instruction[24] _0193_ _0207_ _0240_ i_stall VSS VSS VCC VCC _0391_
+ sky130_fd_sc_hd__a221o_1
X_0730_ _0246_ _0191_ _0261_ i_instruction[2] VSS VSS VCC VCC _0262_ sky130_fd_sc_hd__a22o_1
X_0661_ i_instruction[13] VSS VSS VCC VCC _0198_ sky130_fd_sc_hd__buf_4
X_0592_ o_csr_pc_next[4] i_pc_next[4] _0140_ VSS VSS VCC VCC _0144_ sky130_fd_sc_hd__mux2_1
X_0928_ o_pc[1] i_pc[1] _0151_ VSS VSS VCC VCC _0435_ sky130_fd_sc_hd__mux2_1
X_0859_ _0244_ _0372_ _0373_ _0375_ VSS VSS VCC VCC _0376_ sky130_fd_sc_hd__o22a_1
X_0713_ _0159_ instruction\[6\] _0161_ _0245_ VSS VSS VCC VCC _0022_ sky130_fd_sc_hd__o211a_1
X_0644_ _0177_ _0178_ _0179_ _0180_ _0182_ VSS VSS VCC VCC _0183_ sky130_fd_sc_hd__o41a_2
X_0575_ instruction\[5\] _0064_ _0063_ _0074_ VSS VSS VCC VCC o_reg_write
+ sky130_fd_sc_hd__a31oi_4
X_0627_ _0162_ _0166_ VSS VSS VCC VCC _0167_ sky130_fd_sc_hd__or2_1
X_0558_ _0075_ _0070_ _0099_ o_inst_jal VSS VSS VCC VCC o_op1_src sky130_fd_sc_hd__a31o_2
X_0489_ o_csr_imm[2] _0087_ VSS VSS VCC VCC _0090_ sky130_fd_sc_hd__and2_1
X_0961_ clknet_3_1_0_i_clk _0002_ VSS VSS VCC VCC o_csr_pc_next[3] sky130_fd_sc_hd__dfxtp_2
X_0892_ _0396_ _0403_ _0404_ _0397_ VSS VSS VCC VCC _0405_ sky130_fd_sc_hd__o31a_1
X_0944_ _0443_ VSS VSS VCC VCC _0055_ sky130_fd_sc_hd__clkbuf_1
X_0875_ i_instruction[11] _0189_ _0191_ i_instruction[24] VSS VSS VCC VCC
+ _0390_ sky130_fd_sc_hd__a22o_1
X_0660_ _0163_ i_instruction[8] VSS VSS VCC VCC _0197_ sky130_fd_sc_hd__nand2_2
X_0591_ _0143_ VSS VSS VCC VCC _0002_ sky130_fd_sc_hd__clkbuf_1
X_0927_ o_csr_idx[11] _0349_ _0433_ _0434_ _0161_ VSS VSS VCC VCC _0047_ sky130_fd_sc_hd__o221a_1
X_0858_ _0337_ _0374_ _0196_ VSS VSS VCC VCC _0375_ sky130_fd_sc_hd__o21a_1
X_0789_ _0180_ _0299_ VSS VSS VCC VCC _0314_ sky130_fd_sc_hd__nor2_2
X_0712_ _0240_ _0194_ _0243_ _0244_ _0238_ VSS VSS VCC VCC _0245_ sky130_fd_sc_hd__a221o_1
X_0643_ _0170_ _0181_ _0164_ VSS VSS VCC VCC _0182_ sky130_fd_sc_hd__o21ai_4
X_0574_ _0131_ VSS VSS VCC VCC o_csr_clear sky130_fd_sc_hd__buf_2
X_0626_ _0165_ VSS VSS VCC VCC _0166_ sky130_fd_sc_hd__buf_4
X_0557_ o_csr_imm_sel o_funct3[1] o_funct3[0] _0079_ VSS VSS VCC VCC o_csr_read
+ sky130_fd_sc_hd__o31a_4
X_0488_ _0089_ VSS VSS VCC VCC o_rs1[1] sky130_fd_sc_hd__buf_2
X_0609_ o_csr_pc_next[12] i_pc_next[12] _0151_ VSS VSS VCC VCC _0153_ sky130_fd_sc_hd__mux2_1
X_0960_ clknet_3_7_0_i_clk _0001_ VSS VSS VCC VCC o_csr_pc_next[2] sky130_fd_sc_hd__dfxtp_2
X_0891_ _0246_ _0203_ VSS VSS VCC VCC _0404_ sky130_fd_sc_hd__and2_1
X_0943_ o_pc[8] i_pc[8] _0440_ VSS VSS VCC VCC _0443_ sky130_fd_sc_hd__mux2_1
X_0874_ _0387_ _0388_ _0196_ VSS VSS VCC VCC _0389_ sky130_fd_sc_hd__o21a_1
X_0590_ o_csr_pc_next[3] i_pc_next[3] _0140_ VSS VSS VCC VCC _0143_ sky130_fd_sc_hd__mux2_1
X_0926_ i_instruction[31] _0194_ _0238_ VSS VSS VCC VCC _0434_ sky130_fd_sc_hd__a21o_1
X_0857_ _0212_ _0365_ VSS VSS VCC VCC _0374_ sky130_fd_sc_hd__nor2_1
X_0788_ _0160_ VSS VSS VCC VCC _0313_ sky130_fd_sc_hd__buf_6
X_0711_ _0175_ VSS VSS VCC VCC _0244_ sky130_fd_sc_hd__buf_6
X_0642_ i_instruction[15] VSS VSS VCC VCC _0181_ sky130_fd_sc_hd__buf_6
X_0573_ o_funct3[1] o_funct3[0] _0079_ VSS VSS VCC VCC _0131_ sky130_fd_sc_hd__and3_1
X_0909_ i_instruction[28] _0230_ _0397_ _0419_ _0188_ VSS VSS VCC VCC _0420_
+ sky130_fd_sc_hd__a221o_1
X_0625_ _0164_ VSS VSS VCC VCC _0165_ sky130_fd_sc_hd__buf_4
X_0556_ o_alu_ctrl[3] _0099_ _0118_ VSS VSS VCC VCC o_imm_i[30] sky130_fd_sc_hd__a21o_2
X_0487_ o_csr_imm[1] _0087_ VSS VSS VCC VCC _0089_ sky130_fd_sc_hd__and2_1
X_1039_ o_csr_pc_next[14] VSS VSS VCC VCC o_pc_next[14] sky130_fd_sc_hd__buf_2
X_0608_ _0152_ VSS VSS VCC VCC _0010_ sky130_fd_sc_hd__clkbuf_1
X_0539_ o_csr_imm[0] _0101_ _0120_ VSS VSS VCC VCC o_imm_i[15] sky130_fd_sc_hd__a21o_2
X_0890_ _0222_ _0329_ i_instruction[5] VSS VSS VCC VCC _0403_ sky130_fd_sc_hd__o21a_1
X_0942_ _0442_ VSS VSS VCC VCC _0054_ sky130_fd_sc_hd__clkbuf_1
X_0873_ i_instruction[11] _0203_ _0329_ _0240_ _0337_ VSS VSS VCC VCC _0388_
+ sky130_fd_sc_hd__a221o_1
X_0925_ _0321_ _0423_ _0397_ VSS VSS VCC VCC _0433_ sky130_fd_sc_hd__o21a_1
X_0856_ i_instruction[22] _0193_ _0208_ i_instruction[4] _0188_ vssd1 vssd1 vccd1
+ vccd1 _0373_ sky130_fd_sc_hd__a221o_1
X_0787_ _0159_ o_funct3[1] _0161_ _0312_ VSS VSS VCC VCC _0029_ sky130_fd_sc_hd__o211a_1
X_0710_ _0241_ _0213_ _0242_ _0196_ VSS VSS VCC VCC _0243_ sky130_fd_sc_hd__a2bb2o_1
X_0641_ i_instruction[5] i_instruction[6] _0163_ VSS VSS VCC VCC _0180_ sky130_fd_sc_hd__o21a_1
X_0572_ _0130_ VSS VSS VCC VCC o_csr_set sky130_fd_sc_hd__buf_2
X_0908_ i_instruction[4] _0329_ _0396_ _0418_ VSS VSS VCC VCC _0419_ sky130_fd_sc_hd__a211o_1
X_0839_ i_instruction[15] _0198_ i_ready _0170_ VSS VSS VCC VCC _0358_ sky130_fd_sc_hd__and4bb_4
X_0624_ _0163_ VSS VSS VCC VCC _0164_ sky130_fd_sc_hd__buf_8
X_0555_ o_csr_idx[9] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[29] sky130_fd_sc_hd__a21o_2
X_0486_ _0088_ VSS VSS VCC VCC o_rs1[0] sky130_fd_sc_hd__buf_2
X_1038_ o_csr_pc_next[13] VSS VSS VCC VCC o_pc_next[13] sky130_fd_sc_hd__buf_2
X_0607_ o_csr_pc_next[11] i_pc_next[11] _0151_ VSS VSS VCC VCC _0152_ sky130_fd_sc_hd__mux2_1
X_0538_ o_csr_imm_sel _0101_ _0120_ VSS VSS VCC VCC o_imm_i[14] sky130_fd_sc_hd__a21o_2
X_0469_ _0075_ _0064_ _0076_ VSS VSS VCC VCC _0077_ sky130_fd_sc_hd__and3_1
X_0941_ o_pc[7] i_pc[7] _0440_ VSS VSS VCC VCC _0442_ sky130_fd_sc_hd__mux2_1
X_0872_ _0248_ _0386_ _0358_ _0240_ _0166_ VSS VSS VCC VCC _0387_ sky130_fd_sc_hd__o311a_1
X_0924_ _0349_ o_alu_ctrl[3] _0160_ _0432_ VSS VSS VCC VCC _0046_ sky130_fd_sc_hd__o211a_1
X_0855_ i_instruction[22] _0191_ _0250_ i_instruction[4] _0371_ vssd1 vssd1 vccd1
+ vccd1 _0372_ sky130_fd_sc_hd__a221o_1
X_0786_ _0244_ _0310_ _0311_ _0273_ _0238_ VSS VSS VCC VCC _0312_ sky130_fd_sc_hd__a221o_1
X_0640_ _0163_ i_instruction[12] VSS VSS VCC VCC _0179_ sky130_fd_sc_hd__and2_4
X_0571_ o_funct3[0] _0079_ o_funct3[1] VSS VSS VCC VCC _0130_ sky130_fd_sc_hd__and3b_1
X_0907_ i_instruction[9] _0203_ _0222_ i_instruction[12] VSS VSS VCC VCC _0418_
+ sky130_fd_sc_hd__a22o_1
X_0838_ _0303_ _0295_ VSS VSS VCC VCC _0357_ sky130_fd_sc_hd__nand2_1
X_0769_ _0200_ _0295_ VSS VSS VCC VCC _0296_ sky130_fd_sc_hd__nor2_1
X_0623_ i_ready VSS VSS VCC VCC _0163_ sky130_fd_sc_hd__buf_4
X_0554_ o_csr_idx[8] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[28] sky130_fd_sc_hd__a21o_2
X_0485_ o_csr_imm[0] _0087_ VSS VSS VCC VCC _0088_ sky130_fd_sc_hd__and2_1
X_1037_ o_csr_pc_next[12] VSS VSS VCC VCC o_pc_next[12] sky130_fd_sc_hd__buf_2
X_0606_ _0139_ VSS VSS VCC VCC _0151_ sky130_fd_sc_hd__buf_12
X_0537_ o_funct3[1] _0101_ _0120_ VSS VSS VCC VCC o_imm_i[13] sky130_fd_sc_hd__a21o_2
X_0468_ instruction\[3\] VSS VSS VCC VCC _0076_ sky130_fd_sc_hd__clkinv_2
X_0940_ _0441_ VSS VSS VCC VCC _0053_ sky130_fd_sc_hd__clkbuf_1
X_0871_ _0273_ _0233_ VSS VSS VCC VCC _0386_ sky130_fd_sc_hd__nor2_1
X_0923_ i_instruction[30] _0194_ _0397_ _0431_ _0238_ VSS VSS VCC VCC _0432_
+ sky130_fd_sc_hd__a221o_1
X_0854_ _0181_ _0240_ _0166_ VSS VSS VCC VCC _0371_ sky130_fd_sc_hd__and3b_1
X_0785_ _0175_ _0182_ VSS VSS VCC VCC _0311_ sky130_fd_sc_hd__nor2_2
X_0570_ _0129_ VSS VSS VCC VCC o_csr_write sky130_fd_sc_hd__buf_2
X_0906_ _0168_ _0416_ _0417_ _0216_ VSS VSS VCC VCC _0043_ sky130_fd_sc_hd__o211a_1
X_0837_ i_instruction[2] _0250_ _0355_ _0190_ _0303_ VSS VSS VCC VCC _0356_
+ sky130_fd_sc_hd__a221o_1
X_0768_ _0165_ i_instruction[2] VSS VSS VCC VCC _0295_ sky130_fd_sc_hd__nand2_1
X_0699_ _0164_ _0232_ i_instruction[11] VSS VSS VCC VCC _0233_ sky130_fd_sc_hd__and3_1
X_0622_ i_stall VSS VSS VCC VCC _0162_ sky130_fd_sc_hd__buf_6
X_0553_ o_csr_idx[7] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[27] sky130_fd_sc_hd__a21o_2
X_0484_ _0086_ VSS VSS VCC VCC _0087_ sky130_fd_sc_hd__buf_12
X_1036_ o_csr_pc_next[11] VSS VSS VCC VCC o_pc_next[11] sky130_fd_sc_hd__buf_2
X_0605_ _0150_ VSS VSS VCC VCC _0009_ sky130_fd_sc_hd__clkbuf_1
X_0536_ o_funct3[0] _0101_ _0120_ VSS VSS VCC VCC o_imm_i[12] sky130_fd_sc_hd__a21o_2
X_0467_ instruction\[6\] VSS VSS VCC VCC _0075_ sky130_fd_sc_hd__inv_2
X_1019_ clknet_3_5_0_i_clk _0060_ VSS VSS VCC VCC o_pc[13] sky130_fd_sc_hd__dfxtp_2
X_0519_ _0110_ VSS VSS VCC VCC o_imm_i[5] sky130_fd_sc_hd__buf_2
X_0870_ _0349_ o_csr_idx[3] _0313_ _0385_ VSS VSS VCC VCC _0039_ sky130_fd_sc_hd__o211a_1
X_0999_ clknet_3_0_0_i_clk _0040_ VSS VSS VCC VCC o_csr_idx[4] sky130_fd_sc_hd__dfxtp_4
X_0922_ _0231_ _0429_ _0430_ VSS VSS VCC VCC _0431_ sky130_fd_sc_hd__a21o_1
X_0853_ _0349_ o_csr_idx[1] _0313_ _0370_ VSS VSS VCC VCC _0037_ sky130_fd_sc_hd__o211a_1
X_0784_ _0198_ _0193_ _0207_ _0171_ _0309_ VSS VSS VCC VCC _0310_ sky130_fd_sc_hd__a221o_1
X_0905_ _0157_ o_csr_idx[7] VSS VSS VCC VCC _0417_ sky130_fd_sc_hd__or2_1
X_0836_ _0177_ _0178_ _0253_ _0213_ _0295_ VSS VSS VCC VCC _0355_ sky130_fd_sc_hd__o41ai_1
X_0767_ _0159_ o_rd[4] _0161_ _0294_ VSS VSS VCC VCC _0027_ sky130_fd_sc_hd__o211a_1
X_0698_ i_instruction[10] VSS VSS VCC VCC _0232_ sky130_fd_sc_hd__clkbuf_8
X_0621_ _0160_ VSS VSS VCC VCC _0161_ sky130_fd_sc_hd__buf_6
X_0552_ o_csr_idx[6] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[26] sky130_fd_sc_hd__a21o_2
X_0483_ _0064_ instruction\[3\] _0085_ VSS VSS VCC VCC _0086_ sky130_fd_sc_hd__or3_4
X_1035_ o_csr_pc_next[10] VSS VSS VCC VCC o_pc_next[10] sky130_fd_sc_hd__buf_2
X_0819_ _0171_ _0281_ _0206_ i_instruction[17] VSS VSS VCC VCC _0341_ sky130_fd_sc_hd__a22o_1
X_0604_ o_csr_pc_next[10] i_pc_next[10] _0140_ VSS VSS VCC VCC _0150_ sky130_fd_sc_hd__mux2_1
X_0535_ _0119_ VSS VSS VCC VCC _0120_ sky130_fd_sc_hd__buf_12
X_0466_ instruction\[1\] instruction\[0\] VSS VSS VCC VCC _0074_ sky130_fd_sc_hd__nand2_8
X_1018_ clknet_3_3_0_i_clk _0059_ VSS VSS VCC VCC o_pc[12] sky130_fd_sc_hd__dfxtp_2
X_0518_ o_csr_idx[5] _0086_ VSS VSS VCC VCC _0110_ sky130_fd_sc_hd__and2_1
X_0998_ clknet_3_6_0_i_clk _0039_ VSS VSS VCC VCC o_csr_idx[3] sky130_fd_sc_hd__dfxtp_4
Xclkbuf_3_5_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_5_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0921_ i_instruction[12] _0172_ _0203_ i_instruction[8] _0248_ vssd1 vssd1 vccd1
+ vccd1 _0430_ sky130_fd_sc_hd__a221o_1
X_0852_ _0368_ _0369_ _0168_ VSS VSS VCC VCC _0370_ sky130_fd_sc_hd__a21o_1
X_0783_ _0297_ _0307_ _0308_ _0174_ VSS VSS VCC VCC _0309_ sky130_fd_sc_hd__o31a_1
X_0904_ _0412_ _0414_ _0415_ VSS VSS VCC VCC _0416_ sky130_fd_sc_hd__o21a_1
X_0835_ _0349_ o_csr_imm[4] _0313_ _0354_ VSS VSS VCC VCC _0035_ sky130_fd_sc_hd__o211a_1
X_0766_ _0292_ _0228_ _0293_ _0238_ VSS VSS VCC VCC _0294_ sky130_fd_sc_hd__a31o_1
X_0697_ i_instruction[14] i_instruction[13] i_instruction[15] i_ready vssd1 vssd1
+ vccd1 vccd1 _0231_ sky130_fd_sc_hd__and4bb_4
X_0620_ i_flush VSS VSS VCC VCC _0160_ sky130_fd_sc_hd__clkinv_2
X_0551_ o_csr_idx[5] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[25] sky130_fd_sc_hd__a21o_2
X_0482_ instruction\[2\] VSS VSS VCC VCC _0085_ sky130_fd_sc_hd__inv_2
X_1034_ o_csr_pc_next[9] VSS VSS VCC VCC o_pc_next[9] sky130_fd_sc_hd__buf_2
X_0818_ i_instruction[17] _0230_ _0208_ _0336_ _0339_ VSS VSS VCC VCC _0340_
+ sky130_fd_sc_hd__a221o_1
X_0749_ _0277_ _0278_ _0227_ VSS VSS VCC VCC _0279_ sky130_fd_sc_hd__o21a_1
X_0603_ _0149_ VSS VSS VCC VCC _0008_ sky130_fd_sc_hd__clkbuf_1
X_0534_ _0068_ _0118_ VSS VSS VCC VCC _0119_ sky130_fd_sc_hd__and2b_1
X_0465_ _0072_ _0073_ VSS VSS VCC VCC o_op2_src sky130_fd_sc_hd__nor2_4
X_1017_ clknet_3_5_0_i_clk _0058_ VSS VSS VCC VCC o_pc[11] sky130_fd_sc_hd__dfxtp_2
X_0517_ _0109_ VSS VSS VCC VCC o_imm_i[4] sky130_fd_sc_hd__buf_2
Xclkbuf_3_1_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0997_ clknet_3_2_0_i_clk _0038_ VSS VSS VCC VCC o_csr_idx[2] sky130_fd_sc_hd__dfxtp_4
X_0920_ _0298_ _0292_ _0314_ _0428_ VSS VSS VCC VCC _0429_ sky130_fd_sc_hd__o22a_1
X_0851_ i_instruction[21] _0206_ _0250_ i_instruction[3] _0244_ vssd1 vssd1 vccd1
+ vccd1 _0369_ sky130_fd_sc_hd__a221o_1
X_0782_ _0240_ _0286_ _0231_ i_instruction[11] VSS VSS VCC VCC _0308_ sky130_fd_sc_hd__o211a_1
X_0903_ _0303_ _0177_ _0206_ i_instruction[27] _0175_ VSS VSS VCC VCC _0415_
+ sky130_fd_sc_hd__a221o_1
X_0834_ _0244_ _0352_ _0353_ VSS VSS VCC VCC _0354_ sky130_fd_sc_hd__a21o_1
X_0765_ _0171_ _0188_ _0248_ _0280_ VSS VSS VCC VCC _0293_ sky130_fd_sc_hd__or4_1
X_0696_ _0192_ VSS VSS VCC VCC _0230_ sky130_fd_sc_hd__buf_6
X_0550_ o_csr_idx[4] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[24] sky130_fd_sc_hd__a21o_2
X_0481_ _0084_ VSS VSS VCC VCC o_inst_mret sky130_fd_sc_hd__clkbuf_4
X_1033_ o_csr_pc_next[8] VSS VSS VCC VCC o_pc_next[8] sky130_fd_sc_hd__buf_2
X_0817_ _0321_ _0337_ _0338_ _0282_ VSS VSS VCC VCC _0339_ sky130_fd_sc_hd__o31a_1
X_0748_ i_instruction[9] _0191_ _0250_ _0240_ VSS VSS VCC VCC _0278_ sky130_fd_sc_hd__a22o_1
X_0679_ _0160_ VSS VSS VCC VCC _0216_ sky130_fd_sc_hd__buf_4
X_0602_ o_csr_pc_next[9] i_pc_next[9] _0140_ VSS VSS VCC VCC _0149_ sky130_fd_sc_hd__mux2_1
X_0533_ o_csr_idx[11] _0086_ VSS VSS VCC VCC _0118_ sky130_fd_sc_hd__and2_1
X_0464_ instruction\[6\] _0070_ instruction\[4\] _0063_ o_inst_branch vssd1 vssd1
+ vccd1 vccd1 _0073_ sky130_fd_sc_hd__a41o_1
X_1016_ clknet_3_1_0_i_clk _0057_ VSS VSS VCC VCC o_pc[10] sky130_fd_sc_hd__dfxtp_2
X_0516_ _0087_ _0108_ VSS VSS VCC VCC _0109_ sky130_fd_sc_hd__and2_1
X_0996_ clknet_3_3_0_i_clk _0037_ VSS VSS VCC VCC o_csr_idx[1] sky130_fd_sc_hd__dfxtp_4
X_0850_ i_instruction[21] _0230_ _0367_ _0227_ VSS VSS VCC VCC _0368_ sky130_fd_sc_hd__a211o_1
X_0781_ _0200_ _0211_ VSS VSS VCC VCC _0307_ sky130_fd_sc_hd__nor2_1
X_0979_ clknet_3_0_0_i_clk _0020_ VSS VSS VCC VCC instruction\[4\] sky130_fd_sc_hd__dfxtp_1
X_0902_ i_instruction[27] _0193_ _0208_ _0413_ _0188_ VSS VSS VCC VCC _0414_
+ sky130_fd_sc_hd__a221o_1
X_0833_ i_instruction[19] _0227_ _0206_ _0162_ VSS VSS VCC VCC _0353_ sky130_fd_sc_hd__a31o_1
X_0764_ _0165_ i_instruction[11] VSS VSS VCC VCC _0292_ sky130_fd_sc_hd__and2_2
X_0695_ i_instruction[5] _0171_ _0175_ VSS VSS VCC VCC _0229_ sky130_fd_sc_hd__or3_1
X_0480_ o_csr_idx[2] o_csr_idx[1] _0083_ o_csr_idx[9] VSS VSS VCC VCC _0084_
+ sky130_fd_sc_hd__and4b_1
X_1032_ o_csr_pc_next[7] VSS VSS VCC VCC o_pc_next[7] sky130_fd_sc_hd__buf_2
X_0816_ i_instruction[9] _0220_ _0285_ VSS VSS VCC VCC _0338_ sky130_fd_sc_hd__and3_1
X_0747_ _0267_ _0272_ _0212_ VSS VSS VCC VCC _0277_ sky130_fd_sc_hd__a21oi_1
X_0678_ _0206_ _0208_ _0214_ VSS VSS VCC VCC _0215_ sky130_fd_sc_hd__and3_1
X_0601_ _0148_ VSS VSS VCC VCC _0007_ sky130_fd_sc_hd__clkbuf_1
X_0532_ _0068_ _0116_ _0117_ _0087_ VSS VSS VCC VCC o_imm_i[11] sky130_fd_sc_hd__o211a_2
X_0463_ instruction\[6\] _0071_ VSS VSS VCC VCC _0072_ sky130_fd_sc_hd__nor2_4
X_1015_ clknet_3_6_0_i_clk _0056_ VSS VSS VCC VCC o_pc[9] sky130_fd_sc_hd__dfxtp_2
X_0515_ o_rd[4] o_csr_idx[4] _0096_ VSS VSS VCC VCC _0108_ sky130_fd_sc_hd__mux2_1
X_0995_ clknet_3_3_0_i_clk _0036_ VSS VSS VCC VCC o_csr_idx[0] sky130_fd_sc_hd__dfxtp_4
X_0780_ _0158_ o_funct3[0] _0305_ _0306_ _0216_ VSS VSS VCC VCC _0028_ sky130_fd_sc_hd__o221a_1
X_0978_ clknet_3_0_0_i_clk _0019_ VSS VSS VCC VCC instruction\[3\] sky130_fd_sc_hd__dfxtp_2
X_0901_ i_instruction[3] _0261_ _0250_ i_instruction[8] VSS VSS VCC VCC _0413_
+ sky130_fd_sc_hd__a22o_1
X_0832_ i_instruction[19] _0230_ _0350_ _0351_ VSS VSS VCC VCC _0352_ sky130_fd_sc_hd__a211o_1
X_0763_ _0159_ o_rd[3] _0161_ _0291_ VSS VSS VCC VCC _0026_ sky130_fd_sc_hd__o211a_1
X_0694_ _0227_ _0189_ VSS VSS VCC VCC _0228_ sky130_fd_sc_hd__nand2_1
X_1031_ o_csr_pc_next[6] VSS VSS VCC VCC o_pc_next[6] sky130_fd_sc_hd__buf_2
X_0815_ _0197_ _0178_ _0179_ _0199_ VSS VSS VCC VCC _0337_ sky130_fd_sc_hd__o211a_4
X_0746_ _0158_ o_rd[1] _0266_ _0276_ _0216_ VSS VSS VCC VCC _0024_ sky130_fd_sc_hd__o221a_1
X_0677_ _0209_ _0179_ _0213_ VSS VSS VCC VCC _0214_ sky130_fd_sc_hd__a21oi_2
X_0600_ o_csr_pc_next[8] i_pc_next[8] _0140_ VSS VSS VCC VCC _0148_ sky130_fd_sc_hd__mux2_1
X_0531_ o_csr_idx[0] _0076_ _0065_ VSS VSS VCC VCC _0117_ sky130_fd_sc_hd__or3b_1
X_0462_ _0070_ _0064_ _0063_ VSS VSS VCC VCC _0071_ sky130_fd_sc_hd__or3b_4
X_1014_ clknet_3_5_0_i_clk _0055_ VSS VSS VCC VCC o_pc[8] sky130_fd_sc_hd__dfxtp_2
X_0729_ _0181_ _0219_ VSS VSS VCC VCC _0261_ sky130_fd_sc_hd__nor2_4
X_0514_ _0106_ _0096_ _0107_ VSS VSS VCC VCC o_imm_i[3] sky130_fd_sc_hd__a21oi_4
X_0994_ clknet_3_6_0_i_clk _0035_ VSS VSS VCC VCC o_csr_imm[4] sky130_fd_sc_hd__dfxtp_4
X_0977_ clknet_3_0_0_i_clk _0018_ VSS VSS VCC VCC instruction\[2\] sky130_fd_sc_hd__dfxtp_2
X_0900_ _0396_ _0411_ _0397_ VSS VSS VCC VCC _0412_ sky130_fd_sc_hd__o21a_1
X_0831_ _0189_ _0318_ _0207_ i_instruction[11] _0219_ VSS VSS VCC VCC _0351_
+ sky130_fd_sc_hd__o2111a_1
X_0762_ _0244_ _0288_ _0290_ _0238_ VSS VSS VCC VCC _0291_ sky130_fd_sc_hd__a211o_1
X_0693_ _0188_ VSS VSS VCC VCC _0227_ sky130_fd_sc_hd__buf_6
X_1030_ o_csr_pc_next[5] VSS VSS VCC VCC o_pc_next[5] sky130_fd_sc_hd__buf_2
X_0814_ i_instruction[9] _0191_ _0318_ _0303_ _0281_ VSS VSS VCC VCC _0336_
+ sky130_fd_sc_hd__a32o_1
X_0745_ _0227_ _0269_ _0271_ _0275_ VSS VSS VCC VCC _0276_ sky130_fd_sc_hd__a22o_1
X_0676_ _0210_ _0180_ _0211_ _0212_ VSS VSS VCC VCC _0213_ sky130_fd_sc_hd__or4bb_4
X_0530_ o_rd[0] o_csr_idx[11] _0094_ VSS VSS VCC VCC _0116_ sky130_fd_sc_hd__mux2_1
X_0461_ instruction\[5\] VSS VSS VCC VCC _0070_ sky130_fd_sc_hd__inv_2
X_1013_ clknet_3_3_0_i_clk _0054_ VSS VSS VCC VCC o_pc[7] sky130_fd_sc_hd__dfxtp_2
X_0728_ _0246_ _0230_ _0249_ _0252_ _0259_ VSS VSS VCC VCC _0260_ sky130_fd_sc_hd__a221o_1
X_0659_ _0195_ VSS VSS VCC VCC _0196_ sky130_fd_sc_hd__clkbuf_8
X_0513_ o_rd[3] _0096_ _0087_ VSS VSS VCC VCC _0107_ sky130_fd_sc_hd__o21ai_1
X_0993_ clknet_3_4_0_i_clk _0034_ VSS VSS VCC VCC o_csr_imm[3] sky130_fd_sc_hd__dfxtp_4
X_0976_ clknet_3_2_0_i_clk _0017_ VSS VSS VCC VCC instruction\[1\] sky130_fd_sc_hd__dfxtp_1
X_0830_ _0292_ _0270_ _0321_ _0337_ _0174_ VSS VSS VCC VCC _0350_ sky130_fd_sc_hd__o221a_1
X_0761_ _0183_ _0261_ _0289_ _0188_ VSS VSS VCC VCC _0290_ sky130_fd_sc_hd__o31a_1
X_0692_ _0159_ instruction\[4\] _0161_ _0226_ VSS VSS VCC VCC _0020_ sky130_fd_sc_hd__o211a_1
X_0959_ clknet_3_5_0_i_clk _0000_ VSS VSS VCC VCC o_csr_pc_next[1] sky130_fd_sc_hd__dfxtp_2
X_0813_ _0168_ _0334_ _0335_ _0216_ VSS VSS VCC VCC _0032_ sky130_fd_sc_hd__o211a_1
X_0744_ i_instruction[3] _0250_ _0274_ i_instruction[8] _0248_ VSS VSS VCC VCC
+ _0275_ sky130_fd_sc_hd__a221o_1
X_0675_ _0163_ i_instruction[4] VSS VSS VCC VCC _0212_ sky130_fd_sc_hd__nand2_1
X_0460_ _0069_ VSS VSS VCC VCC o_inst_jal sky130_fd_sc_hd__clkinv_4
X_1012_ clknet_3_0_0_i_clk _0053_ VSS VSS VCC VCC o_pc[6] sky130_fd_sc_hd__dfxtp_2
X_0727_ _0251_ _0257_ _0258_ _0208_ VSS VSS VCC VCC _0259_ sky130_fd_sc_hd__o211a_1
X_0658_ i_instruction[1] _0173_ VSS VSS VCC VCC _0195_ sky130_fd_sc_hd__nor2_4
X_0589_ _0142_ VSS VSS VCC VCC _0001_ sky130_fd_sc_hd__clkbuf_1
X_0512_ o_csr_idx[3] VSS VSS VCC VCC _0106_ sky130_fd_sc_hd__inv_2
X_0992_ clknet_3_4_0_i_clk _0033_ VSS VSS VCC VCC o_csr_imm[2] sky130_fd_sc_hd__dfxtp_4
X_0975_ clknet_3_2_0_i_clk _0016_ VSS VSS VCC VCC instruction\[0\] sky130_fd_sc_hd__dfxtp_1
X_0760_ _0166_ _0232_ _0181_ VSS VSS VCC VCC _0289_ sky130_fd_sc_hd__and3_1
X_0691_ _0218_ _0225_ _0168_ VSS VSS VCC VCC _0226_ sky130_fd_sc_hd__a21o_1
X_0958_ _0450_ VSS VSS VCC VCC _0062_ sky130_fd_sc_hd__clkbuf_1
X_0889_ _0349_ o_csr_idx[5] _0313_ _0402_ VSS VSS VCC VCC _0041_ sky130_fd_sc_hd__o211a_1
X_0812_ _0157_ o_csr_imm[1] VSS VSS VCC VCC _0335_ sky130_fd_sc_hd__or2_1
X_0743_ _0272_ _0273_ VSS VSS VCC VCC _0274_ sky130_fd_sc_hd__nand2_1
X_0674_ _0163_ i_instruction[3] VSS VSS VCC VCC _0211_ sky130_fd_sc_hd__nand2_2
X_1011_ clknet_3_3_0_i_clk _0052_ VSS VSS VCC VCC o_pc[5] sky130_fd_sc_hd__dfxtp_2
X_0726_ _0182_ _0247_ VSS VSS VCC VCC _0258_ sky130_fd_sc_hd__nand2_1
X_0657_ _0188_ _0191_ _0193_ VSS VSS VCC VCC _0194_ sky130_fd_sc_hd__a21o_4
X_0588_ o_csr_pc_next[2] i_pc_next[2] _0140_ VSS VSS VCC VCC _0142_ sky130_fd_sc_hd__mux2_1
X_0511_ _0105_ VSS VSS VCC VCC o_imm_i[2] sky130_fd_sc_hd__buf_2
X_0709_ _0203_ _0222_ VSS VSS VCC VCC _0242_ sky130_fd_sc_hd__or2_1
X_0991_ clknet_3_2_0_i_clk _0032_ VSS VSS VCC VCC o_csr_imm[1] sky130_fd_sc_hd__dfxtp_2
X_0974_ clknet_3_0_0_i_clk _0015_ VSS VSS VCC VCC valid_input sky130_fd_sc_hd__dfxtp_1
X_0690_ _0219_ _0173_ _0221_ _0224_ VSS VSS VCC VCC _0225_ sky130_fd_sc_hd__a31o_1
X_0957_ o_pc[15] i_pc[15] _0440_ VSS VSS VCC VCC _0450_ sky130_fd_sc_hd__mux2_1
X_0888_ _0162_ _0398_ _0400_ _0401_ VSS VSS VCC VCC _0402_ sky130_fd_sc_hd__or4_1
X_0811_ _0328_ _0332_ _0333_ VSS VSS VCC VCC _0334_ sky130_fd_sc_hd__o21a_1
X_0742_ _0198_ _0256_ VSS VSS VCC VCC _0273_ sky130_fd_sc_hd__or2_2
X_0673_ _0163_ i_instruction[2] VSS VSS VCC VCC _0210_ sky130_fd_sc_hd__and2_1
X_1010_ clknet_3_1_0_i_clk _0051_ VSS VSS VCC VCC o_pc[4] sky130_fd_sc_hd__dfxtp_2
X_0725_ _0247_ _0213_ _0254_ _0256_ VSS VSS VCC VCC _0257_ sky130_fd_sc_hd__a211oi_1
X_0656_ _0192_ VSS VSS VCC VCC _0193_ sky130_fd_sc_hd__buf_6
X_0587_ _0141_ VSS VSS VCC VCC _0000_ sky130_fd_sc_hd__clkbuf_1
X_0510_ _0087_ _0104_ VSS VSS VCC VCC _0105_ sky130_fd_sc_hd__and2_1
X_0708_ _0173_ _0190_ VSS VSS VCC VCC _0241_ sky130_fd_sc_hd__nand2_1
X_0639_ i_instruction[7] i_instruction[9] i_instruction[10] i_instruction[11] i_ready
+ VSS VSS VCC VCC _0178_ sky130_fd_sc_hd__o41a_4
X_0990_ clknet_3_4_0_i_clk _0031_ VSS VSS VCC VCC o_csr_imm[0] sky130_fd_sc_hd__dfxtp_4
X_0973_ clknet_3_2_0_i_clk _0014_ VSS VSS VCC VCC o_csr_pc_next[15] sky130_fd_sc_hd__dfxtp_2
X_0956_ _0449_ VSS VSS VCC VCC _0061_ sky130_fd_sc_hd__clkbuf_1
X_0887_ _0171_ _0179_ _0207_ _0193_ i_instruction[25] VSS VSS VCC VCC _0401_
+ sky130_fd_sc_hd__a32o_1
X_0810_ _0171_ _0177_ _0206_ i_instruction[16] _0184_ VSS VSS VCC VCC _0333_
+ sky130_fd_sc_hd__a221o_1
X_0741_ _0181_ _0219_ VSS VSS VCC VCC _0272_ sky130_fd_sc_hd__or2_2
X_0672_ _0177_ _0178_ VSS VSS VCC VCC _0209_ sky130_fd_sc_hd__nor2_1
X_0939_ o_pc[6] i_pc[6] _0440_ VSS VSS VCC VCC _0441_ sky130_fd_sc_hd__mux2_1
X_0724_ _0255_ _0220_ VSS VSS VCC VCC _0256_ sky130_fd_sc_hd__nand2_4
X_0655_ _0173_ _0174_ VSS VSS VCC VCC _0192_ sky130_fd_sc_hd__nor2_2
X_0586_ o_csr_pc_next[1] i_pc_next[1] _0140_ VSS VSS VCC VCC _0141_ sky130_fd_sc_hd__mux2_1
X_0707_ i_instruction[6] VSS VSS VCC VCC _0240_ sky130_fd_sc_hd__buf_4
X_0638_ _0176_ VSS VSS VCC VCC _0177_ sky130_fd_sc_hd__clkbuf_4
X_0569_ o_funct3[1] o_funct3[0] _0079_ VSS VSS VCC VCC _0129_ sky130_fd_sc_hd__and3b_2
X_0972_ clknet_3_7_0_i_clk _0013_ VSS VSS VCC VCC o_csr_pc_next[14] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_3_4_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_4_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0955_ o_pc[14] i_pc[14] _0440_ VSS VSS VCC VCC _0449_ sky130_fd_sc_hd__mux2_1
X_0886_ i_instruction[25] _0256_ _0399_ _0188_ VSS VSS VCC VCC _0400_ sky130_fd_sc_hd__o211a_1
X_0740_ _0177_ _0270_ _0195_ VSS VSS VCC VCC _0271_ sky130_fd_sc_hd__o21a_1
X_0671_ _0207_ VSS VSS VCC VCC _0208_ sky130_fd_sc_hd__buf_4
X_0938_ _0139_ VSS VSS VCC VCC _0440_ sky130_fd_sc_hd__buf_12
X_0869_ _0381_ _0384_ _0168_ VSS VSS VCC VCC _0385_ sky130_fd_sc_hd__a21o_1
X_0723_ _0170_ VSS VSS VCC VCC _0255_ sky130_fd_sc_hd__inv_2
X_0654_ _0190_ VSS VSS VCC VCC _0191_ sky130_fd_sc_hd__buf_4
X_0585_ _0139_ VSS VSS VCC VCC _0140_ sky130_fd_sc_hd__buf_12
X_0706_ _0159_ instruction\[5\] _0161_ _0239_ VSS VSS VCC VCC _0021_ sky130_fd_sc_hd__o211a_1
X_0637_ i_ready i_instruction[8] VSS VSS VCC VCC _0176_ sky130_fd_sc_hd__and2_1
X_0568_ _0128_ VSS VSS VCC VCC o_alu_ctrl[0] sky130_fd_sc_hd__buf_2
X_0499_ _0095_ VSS VSS VCC VCC _0096_ sky130_fd_sc_hd__buf_12
Xclkbuf_3_0_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0971_ clknet_3_0_0_i_clk _0012_ VSS VSS VCC VCC o_csr_pc_next[13] sky130_fd_sc_hd__dfxtp_2
X_0954_ _0448_ VSS VSS VCC VCC _0060_ sky130_fd_sc_hd__clkbuf_1
X_0885_ _0253_ _0256_ VSS VSS VCC VCC _0399_ sky130_fd_sc_hd__nand2_1
X_0670_ i_instruction[0] _0174_ VSS VSS VCC VCC _0207_ sky130_fd_sc_hd__nor2_8
X_0937_ _0439_ VSS VSS VCC VCC _0052_ sky130_fd_sc_hd__clkbuf_1
X_0868_ _0166_ i_instruction[5] _0303_ _0383_ _0175_ VSS VSS VCC VCC _0384_
+ sky130_fd_sc_hd__a311o_1
X_0799_ _0166_ i_instruction[5] _0201_ _0322_ VSS VSS VCC VCC _0323_ sky130_fd_sc_hd__a31o_1
X_0722_ _0209_ _0253_ _0213_ VSS VSS VCC VCC _0254_ sky130_fd_sc_hd__o21ba_1
X_0653_ _0171_ _0189_ VSS VSS VCC VCC _0190_ sky130_fd_sc_hd__nor2_2
X_0584_ i_stall i_flush VSS VSS VCC VCC _0139_ sky130_fd_sc_hd__nor2_4
X_0705_ _0228_ _0229_ _0237_ _0238_ VSS VSS VCC VCC _0239_ sky130_fd_sc_hd__a31o_1
X_0636_ _0173_ _0174_ VSS VSS VCC VCC _0175_ sky130_fd_sc_hd__nand2_4
X_0567_ o_csr_idx[5] o_csr_imm_sel _0072_ VSS VSS VCC VCC _0128_ sky130_fd_sc_hd__and3_1
X_0498_ _0093_ _0094_ VSS VSS VCC VCC _0095_ sky130_fd_sc_hd__and2_1
X_0619_ _0158_ VSS VSS VCC VCC _0159_ sky130_fd_sc_hd__buf_4
X_0970_ clknet_3_7_0_i_clk _0011_ VSS VSS VCC VCC o_csr_pc_next[12] sky130_fd_sc_hd__dfxtp_2
X_0953_ o_pc[13] i_pc[13] _0440_ VSS VSS VCC VCC _0448_ sky130_fd_sc_hd__mux2_1
X_0884_ _0393_ _0396_ _0397_ VSS VSS VCC VCC _0398_ sky130_fd_sc_hd__o21a_1
X_0936_ o_pc[5] i_pc[5] _0151_ VSS VSS VCC VCC _0439_ sky130_fd_sc_hd__mux2_1
X_0867_ _0171_ i_instruction[23] _0220_ _0232_ _0382_ VSS VSS VCC VCC _0383_
+ sky130_fd_sc_hd__o221a_1
X_0798_ _0246_ _0220_ _0285_ _0321_ VSS VSS VCC VCC _0322_ sky130_fd_sc_hd__a31o_1
X_0721_ _0165_ i_instruction[12] VSS VSS VCC VCC _0253_ sky130_fd_sc_hd__nand2_2
X_0652_ _0164_ _0181_ VSS VSS VCC VCC _0189_ sky130_fd_sc_hd__nand2_8
X_0583_ _0138_ VSS VSS VCC VCC o_inst_supported sky130_fd_sc_hd__buf_2
X_0919_ _0232_ _0253_ _0292_ VSS VSS VCC VCC _0428_ sky130_fd_sc_hd__o21ai_1
X_0704_ _0162_ VSS VSS VCC VCC _0238_ sky130_fd_sc_hd__buf_6
X_0635_ _0164_ i_instruction[1] VSS VSS VCC VCC _0174_ sky130_fd_sc_hd__nand2_8
X_0566_ o_alu_ctrl[3] _0124_ _0125_ _0127_ o_inst_branch VSS VSS VCC VCC o_alu_ctrl[2]
+ sky130_fd_sc_hd__a311o_4
X_0497_ instruction\[3\] _0074_ instruction\[2\] _0065_ VSS VSS VCC VCC _0094_
+ sky130_fd_sc_hd__or4b_2
X_0618_ _0157_ VSS VSS VCC VCC _0158_ sky130_fd_sc_hd__buf_4
X_0549_ o_csr_idx[3] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[23] sky130_fd_sc_hd__a21o_2
X_0952_ _0447_ VSS VSS VCC VCC _0059_ sky130_fd_sc_hd__clkbuf_1
X_0883_ _0179_ _0270_ _0195_ VSS VSS VCC VCC _0397_ sky130_fd_sc_hd__o21a_2
X_0935_ _0438_ VSS VSS VCC VCC _0051_ sky130_fd_sc_hd__clkbuf_1
X_0866_ _0182_ VSS VSS VCC VCC _0382_ sky130_fd_sc_hd__inv_2
X_0797_ _0248_ _0297_ VSS VSS VCC VCC _0321_ sky130_fd_sc_hd__or2_4
X_0720_ i_instruction[12] _0250_ _0231_ _0246_ _0251_ VSS VSS VCC VCC _0252_
+ sky130_fd_sc_hd__a221o_1
X_0651_ _0187_ VSS VSS VCC VCC _0188_ sky130_fd_sc_hd__buf_6
X_0582_ _0081_ o_inst_mret _0135_ _0137_ VSS VSS VCC VCC _0138_ sky130_fd_sc_hd__or4b_4
X_0918_ _0349_ o_csr_idx[9] _0313_ _0427_ VSS VSS VCC VCC _0045_ sky130_fd_sc_hd__o211a_1
X_0849_ i_instruction[3] _0272_ _0207_ _0366_ _0196_ VSS VSS VCC VCC _0367_
+ sky130_fd_sc_hd__a32o_1
X_0703_ i_instruction[5] _0230_ _0236_ VSS VSS VCC VCC _0237_ sky130_fd_sc_hd__a21o_1
X_0634_ _0164_ i_instruction[0] VSS VSS VCC VCC _0173_ sky130_fd_sc_hd__nand2_4
X_0565_ o_csr_imm_sel o_funct3[1] _0126_ VSS VSS VCC VCC _0127_ sky130_fd_sc_hd__and3b_1
X_0496_ _0093_ VSS VSS VCC VCC o_inst_store sky130_fd_sc_hd__inv_2
X_0617_ i_stall VSS VSS VCC VCC _0157_ sky130_fd_sc_hd__inv_2
X_0548_ o_csr_idx[2] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[22] sky130_fd_sc_hd__a21o_2
X_0479_ _0080_ VSS VSS VCC VCC _0083_ sky130_fd_sc_hd__inv_2
X_0951_ o_pc[12] i_pc[12] _0440_ VSS VSS VCC VCC _0447_ sky130_fd_sc_hd__mux2_1
X_0882_ _0337_ _0394_ _0395_ VSS VSS VCC VCC _0396_ sky130_fd_sc_hd__or3_2
X_0934_ o_pc[4] i_pc[4] _0151_ VSS VSS VCC VCC _0438_ sky130_fd_sc_hd__mux2_1
X_0865_ _0196_ _0379_ _0380_ _0227_ VSS VSS VCC VCC _0381_ sky130_fd_sc_hd__a211o_1
X_0796_ _0208_ _0258_ _0319_ VSS VSS VCC VCC _0320_ sky130_fd_sc_hd__and3_1
X_0650_ _0173_ _0174_ VSS VSS VCC VCC _0187_ sky130_fd_sc_hd__and2_2
X_0581_ _0067_ _0074_ _0136_ _0094_ valid_input VSS VSS VCC VCC _0137_ sky130_fd_sc_hd__o311a_2
X_0917_ i_instruction[29] _0230_ _0397_ _0424_ _0426_ VSS VSS VCC VCC _0427_
+ sky130_fd_sc_hd__a221o_1
X_0848_ _0211_ _0365_ _0337_ VSS VSS VCC VCC _0366_ sky130_fd_sc_hd__o21bai_1
X_0779_ i_instruction[12] _0227_ _0206_ _0162_ VSS VSS VCC VCC _0306_ sky130_fd_sc_hd__a31o_1
X_0702_ _0181_ _0174_ _0235_ _0173_ VSS VSS VCC VCC _0236_ sky130_fd_sc_hd__o22a_1
X_0633_ _0165_ _0171_ VSS VSS VCC VCC _0172_ sky130_fd_sc_hd__and2_4
X_0564_ o_csr_idx[5] instruction\[6\] _0071_ _0125_ VSS VSS VCC VCC _0126_
+ sky130_fd_sc_hd__o31ai_1
X_0495_ instruction\[5\] _0077_ VSS VSS VCC VCC _0093_ sky130_fd_sc_hd__nand2_2
X_0616_ _0156_ VSS VSS VCC VCC _0014_ sky130_fd_sc_hd__clkbuf_1
X_0547_ o_csr_idx[1] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[21] sky130_fd_sc_hd__a21o_2
X_0478_ _0082_ VSS VSS VCC VCC o_csr_ebreak sky130_fd_sc_hd__buf_2
X_0950_ _0446_ VSS VSS VCC VCC _0058_ sky130_fd_sc_hd__clkbuf_1
X_0881_ _0232_ i_instruction[11] _0179_ _0231_ VSS VSS VCC VCC _0395_ sky130_fd_sc_hd__and4b_1
X_0933_ _0437_ VSS VSS VCC VCC _0050_ sky130_fd_sc_hd__clkbuf_1
X_0864_ i_instruction[23] _0193_ _0207_ i_instruction[5] VSS VSS VCC VCC _0380_
+ sky130_fd_sc_hd__a22o_1
X_0795_ _0246_ _0190_ _0318_ _0303_ VSS VSS VCC VCC _0319_ sky130_fd_sc_hd__a31o_1
X_0580_ o_csr_imm_sel o_funct3[1] o_funct3[0] _0076_ VSS VSS VCC VCC _0136_
+ sky130_fd_sc_hd__o31a_1
X_0916_ _0188_ _0425_ _0162_ VSS VSS VCC VCC _0426_ sky130_fd_sc_hd__a21o_1
X_0847_ _0219_ _0358_ VSS VSS VCC VCC _0365_ sky130_fd_sc_hd__nor2_2
X_0778_ _0302_ _0304_ _0244_ VSS VSS VCC VCC _0305_ sky130_fd_sc_hd__o21a_1
X_0701_ _0200_ _0223_ _0234_ i_instruction[1] VSS VSS VCC VCC _0235_ sky130_fd_sc_hd__a31oi_1
X_0632_ _0170_ VSS VSS VCC VCC _0171_ sky130_fd_sc_hd__buf_6
X_0563_ instruction\[6\] instruction\[5\] _0064_ _0063_ VSS VSS VCC VCC _0125_
+ sky130_fd_sc_hd__or4b_1
X_0494_ _0092_ VSS VSS VCC VCC o_rs1[4] sky130_fd_sc_hd__buf_2
X_0615_ o_csr_pc_next[15] i_pc_next[15] _0151_ VSS VSS VCC VCC _0156_ sky130_fd_sc_hd__mux2_1
X_0546_ o_csr_idx[0] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[20] sky130_fd_sc_hd__a21o_2
X_0477_ o_csr_idx[0] _0081_ VSS VSS VCC VCC _0082_ sky130_fd_sc_hd__and2_4
X_1029_ o_csr_pc_next[4] VSS VSS VCC VCC o_pc_next[4] sky130_fd_sc_hd__buf_2
X_0529_ _0115_ VSS VSS VCC VCC o_imm_i[10] sky130_fd_sc_hd__buf_2
X_0880_ i_instruction[12] _0358_ _0248_ VSS VSS VCC VCC _0394_ sky130_fd_sc_hd__a21o_1
X_0932_ o_pc[3] i_pc[3] _0151_ VSS VSS VCC VCC _0437_ sky130_fd_sc_hd__mux2_1
X_0863_ _0365_ _0378_ _0337_ VSS VSS VCC VCC _0379_ sky130_fd_sc_hd__o21bai_1
X_0794_ _0253_ _0213_ VSS VSS VCC VCC _0318_ sky130_fd_sc_hd__nand2_2
X_0915_ _0303_ _0298_ _0191_ i_instruction[29] VSS VSS VCC VCC _0425_ sky130_fd_sc_hd__a22o_1
X_0846_ _0349_ o_csr_idx[0] _0313_ _0364_ VSS VSS VCC VCC _0036_ sky130_fd_sc_hd__o211a_1
X_0777_ i_instruction[12] _0230_ _0208_ _0303_ VSS VSS VCC VCC _0304_ sky130_fd_sc_hd__a22o_1
X_0700_ _0231_ _0233_ VSS VSS VCC VCC _0234_ sky130_fd_sc_hd__nand2_1
X_0631_ i_instruction[14] VSS VSS VCC VCC _0170_ sky130_fd_sc_hd__clkbuf_8
X_0562_ _0124_ VSS VSS VCC VCC o_alu_ctrl[4] sky130_fd_sc_hd__inv_2
X_0493_ o_csr_imm[4] _0087_ VSS VSS VCC VCC _0092_ sky130_fd_sc_hd__and2_1
X_1045_ o_csr_idx[4] VSS VSS VCC VCC o_rs2[4] sky130_fd_sc_hd__buf_2
X_0829_ _0157_ VSS VSS VCC VCC _0349_ sky130_fd_sc_hd__buf_4
X_0614_ _0155_ VSS VSS VCC VCC _0013_ sky130_fd_sc_hd__clkbuf_1
X_0545_ _0118_ VSS VSS VCC VCC _0122_ sky130_fd_sc_hd__buf_12
X_0476_ o_csr_idx[8] _0080_ VSS VSS VCC VCC _0081_ sky130_fd_sc_hd__nor2_1
X_1028_ o_csr_pc_next[3] VSS VSS VCC VCC o_pc_next[3] sky130_fd_sc_hd__buf_2
X_0528_ o_alu_ctrl[3] _0086_ VSS VSS VCC VCC _0115_ sky130_fd_sc_hd__and2_1
X_0459_ instruction\[2\] _0068_ VSS VSS VCC VCC _0069_ sky130_fd_sc_hd__nand2_1
X_0931_ _0436_ VSS VSS VCC VCC _0049_ sky130_fd_sc_hd__clkbuf_1
X_0862_ _0166_ i_instruction[5] _0234_ VSS VSS VCC VCC _0378_ sky130_fd_sc_hd__a21boi_1
X_0793_ _0159_ o_csr_imm_sel _0313_ _0317_ VSS VSS VCC VCC _0030_ sky130_fd_sc_hd__o211a_1
X_0914_ _0232_ _0203_ _0248_ _0423_ VSS VSS VCC VCC _0424_ sky130_fd_sc_hd__a211o_1
X_0845_ _0362_ _0363_ _0168_ VSS VSS VCC VCC _0364_ sky130_fd_sc_hd__a21o_1
X_0776_ _0182_ VSS VSS VCC VCC _0303_ sky130_fd_sc_hd__buf_6
X_0630_ _0168_ instruction\[0\] VSS VSS VCC VCC _0169_ sky130_fd_sc_hd__nand2_1
X_0561_ o_inst_jal _0077_ _0099_ VSS VSS VCC VCC _0124_ sky130_fd_sc_hd__nor3_4
X_0492_ _0091_ VSS VSS VCC VCC o_rs1[3] sky130_fd_sc_hd__buf_2
X_1044_ o_csr_idx[3] VSS VSS VCC VCC o_rs2[3] sky130_fd_sc_hd__buf_2
X_0828_ _0158_ o_csr_imm[3] _0344_ _0348_ _0216_ VSS VSS VCC VCC _0034_ sky130_fd_sc_hd__o221a_1
X_0759_ _0174_ _0285_ _0287_ _0280_ _0232_ VSS VSS VCC VCC _0288_ sky130_fd_sc_hd__a32o_1
X_0613_ o_csr_pc_next[14] i_pc_next[14] _0151_ VSS VSS VCC VCC _0155_ sky130_fd_sc_hd__mux2_1
X_0544_ _0099_ VSS VSS VCC VCC _0121_ sky130_fd_sc_hd__buf_12
X_0475_ o_csr_imm_sel o_funct3[1] o_funct3[0] _0079_ VSS VSS VCC VCC _0080_
+ sky130_fd_sc_hd__or4b_4
X_1027_ o_csr_pc_next[2] VSS VSS VCC VCC o_pc_next[2] sky130_fd_sc_hd__buf_2
X_0527_ _0114_ VSS VSS VCC VCC o_imm_i[9] sky130_fd_sc_hd__buf_2
X_0458_ instruction\[3\] _0065_ VSS VSS VCC VCC _0068_ sky130_fd_sc_hd__and2_1
X_0930_ o_pc[2] i_pc[2] _0151_ VSS VSS VCC VCC _0436_ sky130_fd_sc_hd__mux2_1
X_0861_ _0168_ _0376_ _0377_ _0216_ VSS VSS VCC VCC _0038_ sky130_fd_sc_hd__o211a_1
X_0792_ _0171_ _0230_ _0316_ _0238_ VSS VSS VCC VCC _0317_ sky130_fd_sc_hd__a211o_1
Xclkbuf_3_7_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_7_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0913_ i_instruction[12] _0172_ _0395_ VSS VSS VCC VCC _0423_ sky130_fd_sc_hd__a21o_1
X_0844_ i_instruction[20] _0206_ _0250_ i_instruction[2] _0244_ vssd1 vssd1 vccd1
+ vccd1 _0363_ sky130_fd_sc_hd__a221o_1
X_0775_ _0296_ _0297_ _0301_ _0174_ VSS VSS VCC VCC _0302_ sky130_fd_sc_hd__o31a_1
X_0560_ _0123_ VSS VSS VCC VCC o_alu_ctrl[1] sky130_fd_sc_hd__buf_2
X_0491_ o_csr_imm[3] _0087_ VSS VSS VCC VCC _0091_ sky130_fd_sc_hd__and2_1
X_1043_ o_csr_idx[2] VSS VSS VCC VCC o_rs2[2] sky130_fd_sc_hd__buf_2
X_0827_ _0208_ _0345_ _0347_ VSS VSS VCC VCC _0348_ sky130_fd_sc_hd__a21o_1
X_0758_ _0286_ _0256_ VSS VSS VCC VCC _0287_ sky130_fd_sc_hd__nand2_1
X_0689_ i_instruction[4] _0192_ _0195_ _0223_ _0187_ VSS VSS VCC VCC _0224_
+ sky130_fd_sc_hd__a221o_1
X_0612_ _0154_ VSS VSS VCC VCC _0012_ sky130_fd_sc_hd__clkbuf_1
X_0543_ o_csr_imm[4] _0101_ _0120_ VSS VSS VCC VCC o_imm_i[19] sky130_fd_sc_hd__a21o_2
X_0474_ _0075_ _0071_ _0074_ VSS VSS VCC VCC _0079_ sky130_fd_sc_hd__nor3_4
X_1026_ o_csr_pc_next[1] VSS VSS VCC VCC o_pc_next[1] sky130_fd_sc_hd__buf_2
X_0526_ o_csr_idx[9] _0086_ VSS VSS VCC VCC _0114_ sky130_fd_sc_hd__and2_1
X_0457_ instruction\[3\] _0067_ VSS VSS VCC VCC o_inst_jalr sky130_fd_sc_hd__nor2_4
X_1009_ clknet_3_5_0_i_clk _0050_ VSS VSS VCC VCC o_pc[3] sky130_fd_sc_hd__dfxtp_2
X_0509_ o_rd[2] o_csr_idx[2] _0096_ VSS VSS VCC VCC _0104_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_3_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_3_3_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0860_ _0157_ o_csr_idx[2] VSS VSS VCC VCC _0377_ sky130_fd_sc_hd__or2_1
X_0791_ _0297_ _0315_ _0196_ VSS VSS VCC VCC _0316_ sky130_fd_sc_hd__o21a_1
X_0989_ clknet_3_1_0_i_clk _0030_ VSS VSS VCC VCC o_csr_imm_sel sky130_fd_sc_hd__dfxtp_4
X_0912_ _0349_ o_csr_idx[8] _0313_ _0422_ VSS VSS VCC VCC _0044_ sky130_fd_sc_hd__o211a_1
X_0843_ _0208_ _0356_ _0357_ _0361_ VSS VSS VCC VCC _0362_ sky130_fd_sc_hd__a31o_1
X_0774_ _0198_ _0250_ _0231_ _0300_ VSS VSS VCC VCC _0301_ sky130_fd_sc_hd__a22o_1
X_0490_ _0090_ VSS VSS VCC VCC o_rs1[2] sky130_fd_sc_hd__buf_2
X_1042_ o_csr_idx[1] VSS VSS VCC VCC o_rs2[1] sky130_fd_sc_hd__buf_2
X_0826_ i_instruction[18] _0193_ _0311_ _0346_ i_stall VSS VSS VCC VCC _0347_
+ sky130_fd_sc_hd__a221o_1
X_0757_ _0165_ _0232_ VSS VSS VCC VCC _0286_ sky130_fd_sc_hd__nand2_1
X_0688_ _0203_ _0222_ VSS VSS VCC VCC _0223_ sky130_fd_sc_hd__nor2_1
X_0611_ o_csr_pc_next[13] i_pc_next[13] _0151_ VSS VSS VCC VCC _0154_ sky130_fd_sc_hd__mux2_1
X_0542_ o_csr_imm[3] _0101_ _0120_ VSS VSS VCC VCC o_imm_i[18] sky130_fd_sc_hd__a21o_2
X_0473_ o_res_src[1] o_res_src[2] VSS VSS VCC VCC o_res_src[0] sky130_fd_sc_hd__nor2_4
X_1025_ o_csr_read VSS VSS VCC VCC o_inst_csr_req sky130_fd_sc_hd__buf_2
X_0809_ i_instruction[16] _0193_ _0271_ _0331_ _0188_ VSS VSS VCC VCC _0332_
+ sky130_fd_sc_hd__a221o_1
X_0525_ _0113_ VSS VSS VCC VCC o_imm_i[8] sky130_fd_sc_hd__buf_2
X_0456_ instruction\[2\] _0065_ VSS VSS VCC VCC _0067_ sky130_fd_sc_hd__nand2_2
X_1008_ clknet_3_0_0_i_clk _0049_ VSS VSS VCC VCC o_pc[2] sky130_fd_sc_hd__dfxtp_2
X_0508_ _0103_ VSS VSS VCC VCC o_imm_i[1] sky130_fd_sc_hd__buf_2
X_0790_ _0200_ _0212_ _0273_ _0314_ VSS VSS VCC VCC _0315_ sky130_fd_sc_hd__o22ai_1
X_0988_ clknet_3_1_0_i_clk _0029_ VSS VSS VCC VCC o_funct3[1] sky130_fd_sc_hd__dfxtp_4
X_0911_ _0420_ _0421_ _0168_ VSS VSS VCC VCC _0422_ sky130_fd_sc_hd__a21o_1
X_0842_ i_instruction[20] _0193_ _0196_ _0360_ _0187_ VSS VSS VCC VCC _0361_
+ sky130_fd_sc_hd__a221o_1
X_0773_ _0165_ i_instruction[5] _0240_ _0299_ VSS VSS VCC VCC _0300_ sky130_fd_sc_hd__a31o_1
X_1041_ o_csr_idx[0] VSS VSS VCC VCC o_rs2[0] sky130_fd_sc_hd__buf_2
X_0825_ i_instruction[18] _0172_ VSS VSS VCC VCC _0346_ sky130_fd_sc_hd__or2_1
X_0756_ _0164_ _0255_ _0198_ VSS VSS VCC VCC _0285_ sky130_fd_sc_hd__nand3_4
X_0687_ _0164_ _0170_ _0181_ VSS VSS VCC VCC _0222_ sky130_fd_sc_hd__and3_2
X_0610_ _0153_ VSS VSS VCC VCC _0011_ sky130_fd_sc_hd__clkbuf_1
X_0541_ o_csr_imm[2] _0101_ _0120_ VSS VSS VCC VCC o_imm_i[17] sky130_fd_sc_hd__a21o_2
X_0472_ _0067_ VSS VSS VCC VCC o_res_src[1] sky130_fd_sc_hd__clkinv_4
X_1024_ o_csr_idx[11] VSS VSS VCC VCC o_imm_i[31] sky130_fd_sc_hd__buf_2
X_0808_ _0166_ _0240_ _0199_ _0329_ _0330_ VSS VSS VCC VCC _0331_ sky130_fd_sc_hd__a311o_1
X_0739_ _0170_ _0181_ _0198_ _0165_ VSS VSS VCC VCC _0270_ sky130_fd_sc_hd__o31a_4
X_0524_ o_csr_idx[8] _0086_ VSS VSS VCC VCC _0113_ sky130_fd_sc_hd__and2_1
X_0455_ _0066_ VSS VSS VCC VCC o_inst_branch sky130_fd_sc_hd__clkbuf_4
X_1007_ clknet_3_7_0_i_clk _0048_ VSS VSS VCC VCC o_pc[1] sky130_fd_sc_hd__dfxtp_2
X_0507_ _0087_ _0102_ VSS VSS VCC VCC _0103_ sky130_fd_sc_hd__and2_1
X_0987_ clknet_3_0_0_i_clk _0028_ VSS VSS VCC VCC o_funct3[0] sky130_fd_sc_hd__dfxtp_4
X_0910_ _0303_ _0281_ _0206_ i_instruction[28] _0244_ VSS VSS VCC VCC _0421_
+ sky130_fd_sc_hd__a221o_1
X_0841_ _0321_ _0337_ _0359_ _0270_ _0210_ VSS VSS VCC VCC _0360_ sky130_fd_sc_hd__o32a_1
X_0772_ i_instruction[11] _0298_ VSS VSS VCC VCC _0299_ sky130_fd_sc_hd__nand2_1
X_1040_ o_csr_pc_next[15] VSS VSS VCC VCC o_pc_next[15] sky130_fd_sc_hd__buf_2
X_0824_ _0232_ _0191_ _0318_ _0303_ _0298_ VSS VSS VCC VCC _0345_ sky130_fd_sc_hd__a32o_1
X_0755_ _0158_ o_rd[2] _0279_ _0284_ _0216_ VSS VSS VCC VCC _0025_ sky130_fd_sc_hd__o221a_1
X_0686_ _0220_ _0214_ VSS VSS VCC VCC _0221_ sky130_fd_sc_hd__nand2_1
X_0540_ o_csr_imm[1] _0101_ _0120_ VSS VSS VCC VCC o_imm_i[16] sky130_fd_sc_hd__a21o_2
X_0471_ _0078_ VSS VSS VCC VCC o_res_src[2] sky130_fd_sc_hd__clkbuf_4
X_1023_ o_csr_imm_sel VSS VSS VCC VCC o_funct3[2] sky130_fd_sc_hd__buf_2
X_0807_ i_instruction[8] _0220_ _0285_ _0321_ VSS VSS VCC VCC _0330_ sky130_fd_sc_hd__a31o_1
X_0738_ i_instruction[8] _0191_ _0261_ i_instruction[3] _0268_ VSS VSS VCC VCC
+ _0269_ sky130_fd_sc_hd__a221o_1
X_0669_ _0191_ VSS VSS VCC VCC _0206_ sky130_fd_sc_hd__buf_4
X_0523_ _0112_ VSS VSS VCC VCC o_imm_i[7] sky130_fd_sc_hd__buf_2
X_0454_ _0063_ _0065_ VSS VSS VCC VCC _0066_ sky130_fd_sc_hd__and2_1
X_1006_ clknet_3_6_0_i_clk _0047_ VSS VSS VCC VCC o_csr_idx[11] sky130_fd_sc_hd__dfxtp_4
X_0506_ o_rd[1] o_csr_idx[1] _0096_ VSS VSS VCC VCC _0102_ sky130_fd_sc_hd__mux2_4
X_0986_ clknet_3_1_0_i_clk _0027_ VSS VSS VCC VCC o_rd[4] sky130_fd_sc_hd__dfxtp_2
X_0840_ _0231_ _0358_ _0210_ VSS VSS VCC VCC _0359_ sky130_fd_sc_hd__o21a_1
X_0771_ _0164_ _0232_ VSS VSS VCC VCC _0298_ sky130_fd_sc_hd__and2_2
X_0969_ clknet_3_3_0_i_clk _0010_ VSS VSS VCC VCC o_csr_pc_next[11] sky130_fd_sc_hd__dfxtp_2
X_0823_ _0298_ _0270_ _0343_ _0196_ VSS VSS VCC VCC _0344_ sky130_fd_sc_hd__o211a_1
X_0754_ i_instruction[9] _0280_ _0282_ _0283_ _0162_ VSS VSS VCC VCC _0284_
+ sky130_fd_sc_hd__a221o_1
X_0685_ _0163_ i_instruction[15] VSS VSS VCC VCC _0220_ sky130_fd_sc_hd__and2_4
X_0470_ _0074_ _0070_ _0077_ VSS VSS VCC VCC _0078_ sky130_fd_sc_hd__and3b_1
X_1022_ o_alu_ctrl[3] VSS VSS VCC VCC o_csr_idx[10] sky130_fd_sc_hd__buf_2
X_0806_ _0197_ _0178_ _0199_ VSS VSS VCC VCC _0329_ sky130_fd_sc_hd__nor3b_4
X_0737_ _0267_ _0211_ VSS VSS VCC VCC _0268_ sky130_fd_sc_hd__nor2_1
X_0668_ i_instruction[2] _0194_ _0196_ _0201_ _0204_ VSS VSS VCC VCC _0205_
+ sky130_fd_sc_hd__a221o_1
X_0599_ _0147_ VSS VSS VCC VCC _0006_ sky130_fd_sc_hd__clkbuf_1
X_0522_ o_csr_idx[7] _0086_ VSS VSS VCC VCC _0112_ sky130_fd_sc_hd__and2_2
X_0453_ instruction\[6\] instruction\[5\] _0064_ VSS VSS VCC VCC _0065_ sky130_fd_sc_hd__and3_1
X_1005_ clknet_3_3_0_i_clk _0046_ VSS VSS VCC VCC o_alu_ctrl[3] sky130_fd_sc_hd__dfxtp_4
X_0505_ _0097_ _0101_ VSS VSS VCC VCC o_imm_i[0] sky130_fd_sc_hd__nor2_4
