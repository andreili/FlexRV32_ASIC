* NGSPICE file created from rv_regs.ext - technology: sky130A

.subckt rv_regs
+ i_clk i_reset_n i_rs_valid i_write
+ i_rs1[0] i_rs1[1] i_rs1[2] i_rs1[3] i_rs1[4] 
+ i_rs2[0] i_rs2[1] i_rs2[2] i_rs2[3] i_rs2[4] 
+ i_rd[0] i_rd[1] i_rd[2] i_rd[3] i_rd[4] 
+ i_data[0] i_data[1] i_data[2] i_data[3] i_data[4] i_data[5] i_data[6] i_data[7] i_data[8] i_data[9] i_data[10] i_data[11] i_data[12] i_data[13] i_data[14] i_data[15] i_data[16] i_data[17] i_data[18] i_data[19] i_data[20] i_data[21] i_data[22] i_data[23] i_data[24] i_data[25] i_data[26] i_data[27] i_data[28] i_data[29] i_data[30] i_data[31] 
+ o_data1[0] o_data1[1] o_data1[2] o_data1[3] o_data1[4] o_data1[5] o_data1[6] o_data1[7] o_data1[8] o_data1[9] o_data1[10] o_data1[11] o_data1[12] o_data1[13] o_data1[14] o_data1[15] o_data1[16] o_data1[17] o_data1[18] o_data1[19] o_data1[20] o_data1[21] o_data1[22] o_data1[23] o_data1[24] o_data1[25] o_data1[26] o_data1[27] o_data1[28] o_data1[29] o_data1[30] o_data1[31] 
+ o_data2[0] o_data2[1] o_data2[2] o_data2[3] o_data2[4] o_data2[5] o_data2[6] o_data2[7] o_data2[8] o_data2[9] o_data2[10] o_data2[11] o_data2[12] o_data2[13] o_data2[14] o_data2[15] o_data2[16] o_data2[17] o_data2[18] o_data2[19] o_data2[20] o_data2[21] o_data2[22] o_data2[23] o_data2[24] o_data2[25] o_data2[26] o_data2[27] o_data2[28] o_data2[29] o_data2[30] o_data2[31] 
+ vccd1 vssd1
X_7963_ _3874_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__clkbuf_1
X_9702_ clknet_leaf_55_i_clk _0846_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6914_ _3311_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__clkbuf_1
X_7894_ _3834_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__clkbuf_1
X_6845_ reg_data\[2\]\[2\] _3133_ _3271_ vssd1 vssd1 vccd1 vccd1 _3274_ sky130_fd_sc_hd__mux2_1
X_9633_ clknet_leaf_7_i_clk _0777_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_9564_ clknet_leaf_76_i_clk _0708_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6776_ i_data[12] vssd1 vssd1 vccd1 vccd1 _3227_ sky130_fd_sc_hd__buf_2
X_8515_ _4178_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__clkbuf_1
X_9495_ clknet_leaf_10_i_clk _0639_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5727_ reg_data\[24\]\[20\] _1847_ _1848_ reg_data\[28\]\[20\] _2312_ vssd1 vssd1
+ vccd1 vccd1 _2313_ sky130_fd_sc_hd__a221o_1
X_8446_ _3923_ reg_data\[17\]\[31\] _4107_ vssd1 vssd1 vccd1 vccd1 _4142_ sky130_fd_sc_hd__mux2_1
X_5658_ _2231_ _2236_ _2241_ _2245_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__or4_1
X_8377_ _4105_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__clkbuf_1
X_4609_ _1162_ _1190_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__and2_4
X_5589_ reg_data\[6\]\[18\] _1951_ _1632_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__and3_1
X_7328_ _3532_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__clkbuf_1
X_7259_ reg_data\[5\]\[2\] _3133_ _3493_ vssd1 vssd1 vccd1 vccd1 _3496_ sky130_fd_sc_hd__mux2_1
X_4960_ reg_data\[3\]\[8\] _1158_ _1567_ _1568_ _1569_ vssd1 vssd1 vccd1 vccd1 _1570_
+ sky130_fd_sc_hd__a2111o_1
X_4891_ reg_data\[26\]\[7\] _1132_ _1134_ reg_data\[29\]\[7\] vssd1 vssd1 vccd1 vccd1
+ _1504_ sky130_fd_sc_hd__a22o_1
X_6630_ i_rd[4] _3121_ _3124_ vssd1 vssd1 vccd1 vccd1 _3125_ sky130_fd_sc_hd__or3_4
X_6561_ r_data2\[2\] _3083_ vssd1 vssd1 vccd1 vccd1 _3086_ sky130_fd_sc_hd__and2_1
X_8300_ _4064_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__clkbuf_1
X_5512_ _2089_ _2094_ _2099_ _2104_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__or4_1
X_9280_ clknet_leaf_70_i_clk _0424_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6492_ r_data1\[2\] _3046_ vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__and2_1
X_8231_ _3913_ reg_data\[14\]\[26\] _4021_ vssd1 vssd1 vccd1 vccd1 _4028_ sky130_fd_sc_hd__mux2_1
X_5443_ reg_data\[6\]\[16\] _1600_ _1716_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__and3_1
X_8162_ _3991_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__clkbuf_1
X_5374_ _1963_ _1967_ _1969_ _1971_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__or4_1
X_7113_ _3266_ reg_data\[8\]\[31\] _3382_ vssd1 vssd1 vccd1 vccd1 _3417_ sky130_fd_sc_hd__mux2_1
X_8093_ _3954_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__clkbuf_1
X_7044_ _3379_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__clkbuf_1
X_8995_ clknet_leaf_64_i_clk _0139_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_7946_ i_data[2] vssd1 vssd1 vccd1 vccd1 _3863_ sky130_fd_sc_hd__clkbuf_4
X_7877_ _3825_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__clkbuf_1
X_9616_ clknet_leaf_31_i_clk _0760_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6828_ i_data[29] vssd1 vssd1 vccd1 vccd1 _3262_ sky130_fd_sc_hd__clkbuf_4
X_9547_ clknet_leaf_27_i_clk _0691_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6759_ _3215_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__clkbuf_1
X_9478_ clknet_leaf_46_i_clk _0622_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8429_ _4133_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_52_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_67_i_clk clknet_3_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5090_ reg_data\[7\]\[10\] _1185_ _1692_ _1694_ _1695_ vssd1 vssd1 vccd1 vccd1 _1696_
+ sky130_fd_sc_hd__a2111o_1
X_8780_ _3917_ reg_data\[29\]\[28\] _4310_ vssd1 vssd1 vccd1 vccd1 _4319_ sky130_fd_sc_hd__mux2_1
X_5992_ reg_data\[16\]\[24\] _2449_ _2450_ reg_data\[9\]\[24\] vssd1 vssd1 vccd1 vccd1
+ _2570_ sky130_fd_sc_hd__a22o_1
X_7800_ _3783_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__clkbuf_1
X_7731_ _3266_ reg_data\[25\]\[31\] _3712_ vssd1 vssd1 vccd1 vccd1 _3747_ sky130_fd_sc_hd__mux2_1
X_4943_ reg_data\[23\]\[8\] _1099_ _1101_ reg_data\[19\]\[8\] vssd1 vssd1 vccd1 vccd1
+ _1554_ sky130_fd_sc_hd__a22o_1
X_7662_ _3710_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__clkbuf_1
X_6613_ r_data2\[27\] _3105_ vssd1 vssd1 vccd1 vccd1 _3113_ sky130_fd_sc_hd__and2_1
X_9401_ clknet_leaf_68_i_clk _0545_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_4874_ reg_data\[3\]\[7\] _1054_ _1484_ _1485_ _1486_ vssd1 vssd1 vccd1 vccd1 _1487_
+ sky130_fd_sc_hd__a2111o_1
X_7593_ _3673_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__clkbuf_1
X_9332_ clknet_leaf_21_i_clk _0476_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6544_ r_data1\[27\] _3068_ vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__and2_1
X_9263_ clknet_leaf_36_i_clk _0407_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6475_ reg_data\[23\]\[1\] _1205_ _1208_ reg_data\[19\]\[1\] vssd1 vssd1 vccd1 vccd1
+ _3035_ sky130_fd_sc_hd__a22o_1
X_8214_ _3896_ reg_data\[14\]\[18\] _4010_ vssd1 vssd1 vccd1 vccd1 _4019_ sky130_fd_sc_hd__mux2_1
X_5426_ reg_data\[1\]\[15\] _1904_ _1905_ reg_data\[15\]\[15\] vssd1 vssd1 vccd1 vccd1
+ _2022_ sky130_fd_sc_hd__a22o_1
X_9194_ clknet_leaf_42_i_clk _0338_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8145_ _3982_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__clkbuf_1
X_5357_ reg_data\[5\]\[14\] _1824_ _1954_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__and3_1
X_5288_ reg_data\[30\]\[13\] _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__and3_1
X_8076_ _3945_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__clkbuf_1
X_7027_ reg_data\[0\]\[23\] _3177_ _3367_ vssd1 vssd1 vccd1 vccd1 _3371_ sky130_fd_sc_hd__mux2_1
X_8978_ clknet_leaf_33_i_clk _0122_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_7929_ _3852_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__clkbuf_1
X_4590_ rs2_mux\[0\] rs2_mux\[1\] vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__nor2_1
X_6260_ reg_data\[1\]\[29\] _2510_ _2511_ reg_data\[15\]\[29\] vssd1 vssd1 vccd1 vccd1
+ _2828_ sky130_fd_sc_hd__a22o_1
X_6191_ reg_data\[18\]\[28\] _2422_ _1167_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__and3_1
X_5211_ reg_data\[17\]\[12\] _1509_ _1275_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__and3_1
X_5142_ reg_data\[6\]\[11\] _1347_ _1632_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__and3_1
X_5073_ _1142_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__clkbuf_4
X_9881_ clknet_leaf_31_i_clk _0951_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_8901_ clknet_leaf_63_i_clk _0045_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8832_ reg_data\[11\]\[20\] i_data[20] _4346_ vssd1 vssd1 vccd1 vccd1 _4347_ sky130_fd_sc_hd__mux2_1
X_5975_ reg_data\[20\]\[24\] _2234_ _1283_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__and3_1
X_8763_ _4287_ vssd1 vssd1 vccd1 vccd1 _4310_ sky130_fd_sc_hd__buf_4
X_7714_ _3738_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__clkbuf_1
X_8694_ _4273_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__clkbuf_1
X_4926_ reg_data\[22\]\[8\] _1536_ _1236_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__and3_1
X_7645_ _3248_ reg_data\[24\]\[22\] _3699_ vssd1 vssd1 vccd1 vccd1 _3702_ sky130_fd_sc_hd__mux2_1
X_4857_ reg_data\[1\]\[6\] _1298_ _1299_ reg_data\[15\]\[6\] vssd1 vssd1 vccd1 vccd1
+ _1471_ sky130_fd_sc_hd__a22o_1
X_7576_ reg_data\[23\]\[22\] _3175_ _3662_ vssd1 vssd1 vccd1 vccd1 _3665_ sky130_fd_sc_hd__mux2_1
X_6527_ r_data1\[19\] _3057_ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__and2_1
X_9315_ clknet_leaf_63_i_clk _0459_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_4788_ reg_data\[20\]\[5\] _1166_ _1180_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__and3_1
X_6458_ reg_data\[22\]\[1\] _1207_ _1151_ vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__and3_1
X_9246_ clknet_leaf_76_i_clk _0390_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6389_ reg_data\[14\]\[0\] _2473_ _1313_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__and3_1
X_5409_ _1142_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__clkbuf_4
X_9177_ clknet_leaf_9_i_clk _0321_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8128_ _3973_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__clkbuf_1
X_8059_ _3936_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__clkbuf_1
X_5760_ reg_data\[22\]\[21\] _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__and3_1
X_5691_ reg_data\[1\]\[20\] _1729_ _1793_ _1794_ reg_data\[15\]\[20\] vssd1 vssd1
+ vccd1 vccd1 _2278_ sky130_fd_sc_hd__a32o_1
X_4711_ reg_data\[27\]\[4\] _1096_ _1327_ _1328_ _1329_ vssd1 vssd1 vccd1 vccd1 _1330_
+ sky130_fd_sc_hd__a2111o_1
X_7430_ _3241_ reg_data\[20\]\[19\] _3576_ vssd1 vssd1 vccd1 vccd1 _3586_ sky130_fd_sc_hd__mux2_1
X_4642_ reg_data\[1\]\[3\] _1022_ _1109_ _1111_ reg_data\[15\]\[3\] vssd1 vssd1 vccd1
+ vccd1 _1263_ sky130_fd_sc_hd__a32o_1
X_7361_ _3549_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__clkbuf_1
X_4573_ reg_data\[7\]\[2\] _1185_ _1188_ _1192_ _1194_ vssd1 vssd1 vccd1 vccd1 _1195_
+ sky130_fd_sc_hd__a2111o_1
X_9100_ clknet_leaf_27_i_clk _0244_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6312_ reg_data\[23\]\[30\] _2440_ _2441_ reg_data\[19\]\[30\] vssd1 vssd1 vccd1
+ vccd1 _2878_ sky130_fd_sc_hd__a22o_1
X_7292_ reg_data\[5\]\[18\] _3166_ _3504_ vssd1 vssd1 vccd1 vccd1 _3513_ sky130_fd_sc_hd__mux2_1
X_6243_ reg_data\[17\]\[29\] _1162_ _1148_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__and3_1
X_9031_ clknet_leaf_52_i_clk _0175_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6174_ reg_data\[13\]\[28\] _2214_ _1087_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__and3_1
X_5125_ reg_data\[1\]\[11\] _1729_ _1109_ _1111_ reg_data\[15\]\[11\] vssd1 vssd1
+ vccd1 vccd1 _1730_ sky130_fd_sc_hd__a32o_1
X_5056_ reg_data\[5\]\[10\] _1490_ _1250_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__and3_1
X_9864_ clknet_leaf_71_i_clk _0934_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_9795_ clknet_leaf_55_i_clk rdata1\[11\] vssd1 vssd1 vccd1 vccd1 r_data1\[11\] sky130_fd_sc_hd__dfxtp_1
X_8815_ reg_data\[11\]\[12\] i_data[12] _4335_ vssd1 vssd1 vccd1 vccd1 _4338_ sky130_fd_sc_hd__mux2_1
X_5958_ _2522_ _2527_ _2532_ _2536_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__or4_1
X_8746_ _4301_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__clkbuf_1
X_4909_ reg_data\[0\]\[7\] _1174_ _1518_ _1519_ _1520_ vssd1 vssd1 vccd1 vccd1 _1521_
+ sky130_fd_sc_hd__a2111o_1
X_5889_ reg_data\[4\]\[23\] _2325_ _2469_ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__and3_1
X_8677_ reg_data\[19\]\[11\] _3152_ _4263_ vssd1 vssd1 vccd1 vccd1 _4265_ sky130_fd_sc_hd__mux2_1
X_7628_ _3231_ reg_data\[24\]\[14\] _3688_ vssd1 vssd1 vccd1 vccd1 _3693_ sky130_fd_sc_hd__mux2_1
X_7559_ reg_data\[23\]\[14\] _3158_ _3651_ vssd1 vssd1 vccd1 vccd1 _3656_ sky130_fd_sc_hd__mux2_1
X_9229_ clknet_leaf_28_i_clk _0373_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6930_ _3319_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__clkbuf_1
X_6861_ _3270_ vssd1 vssd1 vccd1 vccd1 _3282_ sky130_fd_sc_hd__buf_4
X_5812_ reg_data\[23\]\[22\] _2393_ _2394_ reg_data\[19\]\[22\] vssd1 vssd1 vccd1
+ vccd1 _2395_ sky130_fd_sc_hd__a22o_1
X_9580_ clknet_leaf_40_i_clk _0724_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8600_ _3873_ reg_data\[12\]\[7\] _4216_ vssd1 vssd1 vccd1 vccd1 _4224_ sky130_fd_sc_hd__mux2_1
X_6792_ _3237_ reg_data\[22\]\[17\] _3223_ vssd1 vssd1 vccd1 vccd1 _3238_ sky130_fd_sc_hd__mux2_1
X_5743_ reg_data\[0\]\[21\] _1775_ _2324_ _2326_ _2327_ vssd1 vssd1 vccd1 vccd1 _2328_
+ sky130_fd_sc_hd__a2111o_1
X_8531_ _4187_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__clkbuf_1
X_5674_ _1038_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__clkbuf_4
X_8462_ _3871_ reg_data\[18\]\[6\] _4144_ vssd1 vssd1 vccd1 vccd1 _4151_ sky130_fd_sc_hd__mux2_1
X_7413_ _3577_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__clkbuf_1
X_4625_ reg_data\[3\]\[3\] _1054_ _1243_ _1244_ _1245_ vssd1 vssd1 vccd1 vccd1 _1246_
+ sky130_fd_sc_hd__a2111o_1
X_8393_ _4114_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__clkbuf_1
X_4556_ reg_data\[6\]\[2\] _1177_ _1152_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__and3_1
X_7344_ reg_data\[3\]\[10\] _3149_ _3540_ vssd1 vssd1 vccd1 vccd1 _3541_ sky130_fd_sc_hd__mux2_1
X_4487_ _1020_ rs1_mux\[2\] rs1_mux\[3\] _1052_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__and4_4
X_7275_ _3492_ vssd1 vssd1 vccd1 vccd1 _3504_ sky130_fd_sc_hd__clkbuf_8
X_6226_ reg_data\[14\]\[29\] _2473_ _1313_ vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__and3_1
X_9014_ clknet_leaf_16_i_clk _0158_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6157_ reg_data\[24\]\[27\] _2453_ _2454_ reg_data\[28\]\[27\] _2728_ vssd1 vssd1
+ vccd1 vccd1 _2729_ sky130_fd_sc_hd__a221o_1
X_5108_ reg_data\[30\]\[11\] _1312_ _1313_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__and3_1
X_6088_ reg_data\[5\]\[26\] _1175_ _1273_ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__and3_1
X_9916_ clknet_leaf_32_i_clk _0986_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_5039_ reg_data\[8\]\[9\] _1214_ _1217_ reg_data\[10\]\[9\] _1646_ vssd1 vssd1 vccd1
+ vccd1 _1647_ sky130_fd_sc_hd__a221o_1
X_9847_ clknet_leaf_38_i_clk rdata2\[31\] vssd1 vssd1 vccd1 vccd1 r_data2\[31\] sky130_fd_sc_hd__dfxtp_1
X_9778_ clknet_leaf_37_i_clk _0922_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_8729_ _4292_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__clkbuf_1
X_4410_ _1033_ vssd1 vssd1 vccd1 vccd1 rs1_mux\[3\] sky130_fd_sc_hd__inv_2
X_5390_ reg_data\[14\]\[15\] _1986_ _1090_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__and3_1
X_7060_ _3389_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__clkbuf_1
X_6011_ reg_data\[12\]\[25\] _1082_ _2271_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__and3_1
X_7962_ _3873_ reg_data\[9\]\[7\] _3859_ vssd1 vssd1 vccd1 vccd1 _3874_ sky130_fd_sc_hd__mux2_1
X_9701_ clknet_leaf_57_i_clk _0845_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6913_ _3204_ reg_data\[10\]\[1\] _3309_ vssd1 vssd1 vccd1 vccd1 _3311_ sky130_fd_sc_hd__mux2_1
X_7893_ _3222_ reg_data\[28\]\[10\] _3833_ vssd1 vssd1 vccd1 vccd1 _3834_ sky130_fd_sc_hd__mux2_1
X_9632_ clknet_leaf_7_i_clk _0776_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6844_ _3273_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__clkbuf_1
X_9563_ clknet_leaf_76_i_clk _0707_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6775_ _3226_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__clkbuf_1
X_9494_ clknet_leaf_15_i_clk _0638_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_8514_ _3923_ reg_data\[18\]\[31\] _4143_ vssd1 vssd1 vccd1 vccd1 _4178_ sky130_fd_sc_hd__mux2_1
X_5726_ reg_data\[26\]\[20\] _1849_ _1850_ reg_data\[29\]\[20\] vssd1 vssd1 vccd1
+ vccd1 _2312_ sky130_fd_sc_hd__a22o_1
X_8445_ _4141_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__clkbuf_1
X_5657_ reg_data\[7\]\[19\] _1827_ _2242_ _2243_ _2244_ vssd1 vssd1 vccd1 vccd1 _2245_
+ sky130_fd_sc_hd__a2111o_1
X_8376_ _3921_ reg_data\[16\]\[30\] _4071_ vssd1 vssd1 vccd1 vccd1 _4105_ sky130_fd_sc_hd__mux2_1
X_5588_ reg_data\[3\]\[18\] _1815_ _2175_ _2176_ _2177_ vssd1 vssd1 vccd1 vccd1 _2178_
+ sky130_fd_sc_hd__a2111o_1
X_4608_ _1229_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__clkbuf_4
X_7327_ reg_data\[3\]\[2\] _3133_ _3529_ vssd1 vssd1 vccd1 vccd1 _3532_ sky130_fd_sc_hd__mux2_1
X_4539_ reg_data\[20\]\[2\] _1159_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__and3_1
X_7258_ _3495_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__clkbuf_1
X_6209_ reg_data\[8\]\[28\] _2447_ _2448_ reg_data\[10\]\[28\] _2778_ vssd1 vssd1
+ vccd1 vccd1 _2779_ sky130_fd_sc_hd__a221o_1
X_7189_ _3458_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__clkbuf_1
X_4890_ reg_data\[8\]\[7\] _1116_ _1119_ reg_data\[10\]\[7\] _1502_ vssd1 vssd1 vccd1
+ vccd1 _1503_ sky130_fd_sc_hd__a221o_1
X_6560_ _3085_ vssd1 vssd1 vccd1 vccd1 o_data2[1] sky130_fd_sc_hd__buf_2
X_5511_ reg_data\[7\]\[17\] _1780_ _2100_ _2101_ _2103_ vssd1 vssd1 vccd1 vccd1 _2104_
+ sky130_fd_sc_hd__a2111o_1
X_6491_ _3048_ vssd1 vssd1 vccd1 vccd1 o_data1[1] sky130_fd_sc_hd__buf_2
X_8230_ _4027_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__clkbuf_1
X_5442_ reg_data\[3\]\[16\] _1770_ _2033_ _2034_ _2036_ vssd1 vssd1 vccd1 vccd1 _2037_
+ sky130_fd_sc_hd__a2111o_1
X_8161_ _3911_ reg_data\[13\]\[25\] _3985_ vssd1 vssd1 vccd1 vccd1 _3991_ sky130_fd_sc_hd__mux2_1
X_5373_ reg_data\[24\]\[14\] _1847_ _1848_ reg_data\[28\]\[14\] _1970_ vssd1 vssd1
+ vccd1 vccd1 _1971_ sky130_fd_sc_hd__a221o_1
X_8092_ _3911_ reg_data\[30\]\[25\] _3948_ vssd1 vssd1 vccd1 vccd1 _3954_ sky130_fd_sc_hd__mux2_1
X_7112_ _3416_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
X_7043_ reg_data\[0\]\[31\] _3193_ _3344_ vssd1 vssd1 vccd1 vccd1 _3379_ sky130_fd_sc_hd__mux2_1
X_8994_ clknet_leaf_66_i_clk _0138_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_7945_ _3862_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__clkbuf_1
X_7876_ _3206_ reg_data\[28\]\[2\] _3822_ vssd1 vssd1 vccd1 vccd1 _3825_ sky130_fd_sc_hd__mux2_1
X_6827_ _3261_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__clkbuf_1
X_9615_ clknet_leaf_32_i_clk _0759_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_9546_ clknet_leaf_26_i_clk _0690_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6758_ _3214_ reg_data\[22\]\[6\] _3202_ vssd1 vssd1 vccd1 vccd1 _3215_ sky130_fd_sc_hd__mux2_1
X_5709_ reg_data\[6\]\[20\] _1951_ _2237_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__and3_1
X_6689_ i_data[18] vssd1 vssd1 vccd1 vccd1 _3166_ sky130_fd_sc_hd__clkbuf_4
X_9477_ clknet_leaf_65_i_clk _0621_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8428_ _3905_ reg_data\[17\]\[22\] _4130_ vssd1 vssd1 vccd1 vccd1 _4133_ sky130_fd_sc_hd__mux2_1
X_8359_ _4096_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__clkbuf_1
X_5991_ reg_data\[27\]\[24\] _2439_ _2566_ _2567_ _2568_ vssd1 vssd1 vccd1 vccd1 _2569_
+ sky130_fd_sc_hd__a2111o_1
X_7730_ _3746_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__clkbuf_1
X_4942_ _1540_ _1544_ _1548_ _1552_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__or4_1
X_7661_ _3264_ reg_data\[24\]\[30\] _3676_ vssd1 vssd1 vccd1 vccd1 _3710_ sky130_fd_sc_hd__mux2_1
X_6612_ _3112_ vssd1 vssd1 vccd1 vccd1 o_data2[26] sky130_fd_sc_hd__buf_2
X_9400_ clknet_leaf_61_i_clk _0544_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_4873_ reg_data\[20\]\[7\] _1062_ _1315_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__and3_1
X_7592_ reg_data\[23\]\[30\] _3191_ _3639_ vssd1 vssd1 vccd1 vccd1 _3673_ sky130_fd_sc_hd__mux2_1
X_9331_ clknet_leaf_21_i_clk _0475_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6543_ _3075_ vssd1 vssd1 vccd1 vccd1 o_data1[26] sky130_fd_sc_hd__buf_2
X_9262_ clknet_leaf_39_i_clk _0406_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6474_ _3021_ _3025_ _3029_ _3033_ vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__or4_2
X_8213_ _4018_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__clkbuf_1
X_5425_ reg_data\[2\]\[15\] _1837_ _1901_ _1902_ reg_data\[11\]\[15\] vssd1 vssd1
+ vccd1 vccd1 _2021_ sky130_fd_sc_hd__a32o_1
X_9193_ clknet_leaf_41_i_clk _0337_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_5356_ _1144_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__clkbuf_4
X_8144_ _3894_ reg_data\[13\]\[17\] _3974_ vssd1 vssd1 vccd1 vccd1 _3982_ sky130_fd_sc_hd__mux2_1
X_5287_ reg_data\[18\]\[13\] _1816_ _1513_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__and3_1
X_8075_ _3894_ reg_data\[30\]\[17\] _3937_ vssd1 vssd1 vccd1 vccd1 _3945_ sky130_fd_sc_hd__mux2_1
X_7026_ _3370_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__clkbuf_1
X_8977_ clknet_leaf_31_i_clk _0121_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_7928_ _3258_ reg_data\[28\]\[27\] _3844_ vssd1 vssd1 vccd1 vccd1 _3852_ sky130_fd_sc_hd__mux2_1
X_7859_ _3258_ reg_data\[27\]\[27\] _3807_ vssd1 vssd1 vccd1 vccd1 _3815_ sky130_fd_sc_hd__mux2_1
X_9529_ clknet_leaf_12_i_clk _0673_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_5210_ reg_data\[21\]\[12\] _1272_ _1273_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__and3_1
X_6190_ reg_data\[25\]\[28\] _2416_ _2757_ _2758_ _2759_ vssd1 vssd1 vccd1 vccd1 _2760_
+ sky130_fd_sc_hd__a2111o_1
X_5141_ reg_data\[3\]\[11\] _1158_ _1741_ _1742_ _1744_ vssd1 vssd1 vccd1 vccd1 _1745_
+ sky130_fd_sc_hd__a2111o_1
X_5072_ _1678_ vssd1 vssd1 vccd1 vccd1 rdata1\[10\] sky130_fd_sc_hd__clkbuf_1
X_8900_ clknet_leaf_47_i_clk _0044_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_9880_ clknet_leaf_38_i_clk _0950_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_8831_ _4323_ vssd1 vssd1 vccd1 vccd1 _4346_ sky130_fd_sc_hd__buf_4
X_8762_ _4309_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__clkbuf_1
X_5974_ reg_data\[30\]\[24\] _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__and3_1
X_7713_ _3248_ reg_data\[25\]\[22\] _3735_ vssd1 vssd1 vccd1 vccd1 _3738_ sky130_fd_sc_hd__mux2_1
X_8693_ reg_data\[19\]\[19\] _3168_ _4263_ vssd1 vssd1 vccd1 vccd1 _4273_ sky130_fd_sc_hd__mux2_1
X_4925_ _1038_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__clkbuf_4
X_4856_ reg_data\[2\]\[6\] _1002_ _1295_ _1296_ reg_data\[11\]\[6\] vssd1 vssd1 vccd1
+ vccd1 _1470_ sky130_fd_sc_hd__a32o_1
X_7644_ _3701_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__clkbuf_1
X_7575_ _3664_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__clkbuf_1
X_6526_ _3066_ vssd1 vssd1 vccd1 vccd1 o_data1[18] sky130_fd_sc_hd__buf_2
X_9314_ clknet_leaf_64_i_clk _0458_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_51_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4787_ reg_data\[30\]\[5\] _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__and3_1
X_6457_ _3017_ vssd1 vssd1 vccd1 vccd1 rdata1\[1\] sky130_fd_sc_hd__dlymetal6s2s_1
X_9245_ clknet_leaf_0_i_clk _0389_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6388_ reg_data\[0\]\[0\] _1069_ _2948_ _2949_ _2950_ vssd1 vssd1 vccd1 vccd1 _2951_
+ sky130_fd_sc_hd__a2111o_1
X_9176_ clknet_leaf_10_i_clk _0320_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_5408_ reg_data\[18\]\[15\] _1816_ _1513_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__and3_1
X_5339_ reg_data\[8\]\[14\] _1797_ _1798_ reg_data\[10\]\[14\] _1937_ vssd1 vssd1
+ vccd1 vccd1 _1938_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_66_i_clk clknet_3_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_8127_ _3877_ reg_data\[13\]\[9\] _3963_ vssd1 vssd1 vccd1 vccd1 _3973_ sky130_fd_sc_hd__mux2_1
X_8058_ _3877_ reg_data\[30\]\[9\] _3926_ vssd1 vssd1 vccd1 vccd1 _3936_ sky130_fd_sc_hd__mux2_1
X_7009_ _3361_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_19_i_clk clknet_3_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4710_ reg_data\[1\]\[4\] _1022_ _1109_ _1111_ reg_data\[15\]\[4\] vssd1 vssd1 vccd1
+ vccd1 _1329_ sky130_fd_sc_hd__a32o_1
X_5690_ reg_data\[2\]\[20\] _2219_ _1790_ _1791_ reg_data\[11\]\[20\] vssd1 vssd1
+ vccd1 vccd1 _2277_ sky130_fd_sc_hd__a32o_1
X_4641_ reg_data\[2\]\[3\] _1103_ _1104_ _1106_ reg_data\[11\]\[3\] vssd1 vssd1 vccd1
+ vccd1 _1262_ sky130_fd_sc_hd__a32o_1
X_7360_ reg_data\[3\]\[18\] _3166_ _3540_ vssd1 vssd1 vccd1 vccd1 _3549_ sky130_fd_sc_hd__mux2_1
X_4572_ reg_data\[14\]\[2\] _1001_ _1193_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__and3_1
X_6311_ _2864_ _2868_ _2872_ _2876_ vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__or4_4
X_7291_ _3512_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__clkbuf_1
X_6242_ reg_data\[21\]\[29\] _2489_ _1943_ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__and3_1
X_9030_ clknet_leaf_51_i_clk _0174_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6173_ reg_data\[12\]\[28\] _1082_ _2271_ vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__and3_1
X_5124_ _1021_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__buf_4
X_5055_ reg_data\[4\]\[10\] _1074_ _1248_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__and3_1
X_9863_ clknet_leaf_70_i_clk _0933_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_8814_ _4337_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__clkbuf_1
X_9794_ clknet_leaf_54_i_clk rdata1\[10\] vssd1 vssd1 vccd1 vccd1 r_data1\[10\] sky130_fd_sc_hd__dfxtp_1
X_5957_ reg_data\[7\]\[24\] _2386_ _2533_ _2534_ _2535_ vssd1 vssd1 vccd1 vccd1 _2536_
+ sky130_fd_sc_hd__a2111o_1
X_8745_ _3882_ reg_data\[29\]\[11\] _4299_ vssd1 vssd1 vccd1 vccd1 _4301_ sky130_fd_sc_hd__mux2_1
X_8676_ _4264_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__clkbuf_1
X_4908_ reg_data\[5\]\[7\] _1179_ _1285_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__and3_1
X_5888_ _1059_ vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__buf_2
X_7627_ _3692_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__clkbuf_1
X_4839_ reg_data\[17\]\[6\] _1150_ _1275_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__and3_1
X_7558_ _3655_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__clkbuf_1
X_6509_ r_data1\[10\] _3057_ vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__and2_1
X_7489_ _3618_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__clkbuf_1
X_9228_ clknet_leaf_28_i_clk _0372_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_9159_ clknet_leaf_46_i_clk _0303_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6860_ _3281_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__clkbuf_1
X_5811_ _1100_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__buf_2
X_6791_ i_data[17] vssd1 vssd1 vccd1 vccd1 _3237_ sky130_fd_sc_hd__buf_2
X_5742_ reg_data\[5\]\[21\] _2097_ _1925_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__and3_1
X_8530_ reg_data\[1\]\[6\] _3141_ _4180_ vssd1 vssd1 vccd1 vccd1 _4187_ sky130_fd_sc_hd__mux2_1
X_5673_ reg_data\[25\]\[20\] _1764_ _2257_ _2258_ _2259_ vssd1 vssd1 vccd1 vccd1 _2260_
+ sky130_fd_sc_hd__a2111o_1
X_8461_ _4150_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__clkbuf_1
X_7412_ _3222_ reg_data\[20\]\[10\] _3576_ vssd1 vssd1 vccd1 vccd1 _3577_ sky130_fd_sc_hd__mux2_1
X_8392_ _3869_ reg_data\[17\]\[5\] _4108_ vssd1 vssd1 vccd1 vccd1 _4114_ sky130_fd_sc_hd__mux2_1
X_4624_ reg_data\[30\]\[3\] _1062_ _1090_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__and3_1
X_4555_ _1171_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__buf_2
X_7343_ _3528_ vssd1 vssd1 vccd1 vccd1 _3540_ sky130_fd_sc_hd__buf_4
X_9013_ clknet_leaf_16_i_clk _0157_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_4486_ _1108_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__buf_4
X_7274_ _3503_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__clkbuf_1
X_6225_ reg_data\[0\]\[29\] _2381_ _2791_ _2792_ _2793_ vssd1 vssd1 vccd1 vccd1 _2794_
+ sky130_fd_sc_hd__a2111o_1
X_6156_ reg_data\[26\]\[27\] _2455_ _2456_ reg_data\[29\]\[27\] vssd1 vssd1 vccd1
+ vccd1 _2728_ sky130_fd_sc_hd__a22o_1
X_5107_ reg_data\[18\]\[11\] _1656_ _1483_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__and3_1
X_6087_ reg_data\[6\]\[26\] _2555_ _2237_ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__and3_1
X_9915_ clknet_leaf_32_i_clk _0985_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_5038_ reg_data\[16\]\[9\] _1219_ _1221_ reg_data\[9\]\[9\] vssd1 vssd1 vccd1 vccd1
+ _1646_ sky130_fd_sc_hd__a22o_1
X_9846_ clknet_leaf_39_i_clk rdata2\[30\] vssd1 vssd1 vccd1 vccd1 r_data2\[30\] sky130_fd_sc_hd__dfxtp_1
X_9777_ clknet_leaf_35_i_clk _0921_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_8728_ _3865_ reg_data\[29\]\[3\] _4288_ vssd1 vssd1 vccd1 vccd1 _4292_ sky130_fd_sc_hd__mux2_1
X_6989_ reg_data\[0\]\[5\] _3139_ _3345_ vssd1 vssd1 vccd1 vccd1 _3351_ sky130_fd_sc_hd__mux2_1
X_8659_ _4255_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__clkbuf_1
X_6010_ reg_data\[14\]\[25\] _2473_ _2156_ vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__and3_1
X_7961_ i_data[7] vssd1 vssd1 vccd1 vccd1 _3873_ sky130_fd_sc_hd__clkbuf_4
X_6912_ _3310_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__clkbuf_1
X_9700_ clknet_leaf_60_i_clk _0844_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_7892_ _3821_ vssd1 vssd1 vccd1 vccd1 _3833_ sky130_fd_sc_hd__buf_4
X_6843_ reg_data\[2\]\[1\] _3131_ _3271_ vssd1 vssd1 vccd1 vccd1 _3273_ sky130_fd_sc_hd__mux2_1
X_9631_ clknet_leaf_7_i_clk _0775_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_9562_ clknet_leaf_1_i_clk _0706_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6774_ _3225_ reg_data\[22\]\[11\] _3223_ vssd1 vssd1 vccd1 vccd1 _3226_ sky130_fd_sc_hd__mux2_1
X_9493_ clknet_leaf_15_i_clk _0637_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_8513_ _4177_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__clkbuf_1
X_5725_ reg_data\[8\]\[20\] _1841_ _1842_ reg_data\[10\]\[20\] _2310_ vssd1 vssd1
+ vccd1 vccd1 _2311_ sky130_fd_sc_hd__a221o_1
X_8444_ _3921_ reg_data\[17\]\[30\] _4107_ vssd1 vssd1 vccd1 vccd1 _4141_ sky130_fd_sc_hd__mux2_1
X_5656_ reg_data\[13\]\[19\] _1960_ _1191_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__and3_1
X_4607_ _1207_ _1215_ _1197_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__and3_4
X_8375_ _4104_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__clkbuf_1
X_5587_ reg_data\[30\]\[18\] _1629_ _1344_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__and3_1
X_4538_ _0993_ _1006_ rs2_mux\[2\] _1013_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__and4_4
X_7326_ _3531_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__clkbuf_1
X_7257_ reg_data\[5\]\[1\] _3131_ _3493_ vssd1 vssd1 vccd1 vccd1 _3495_ sky130_fd_sc_hd__mux2_1
X_4469_ reg_data\[7\]\[2\] _1081_ _1084_ _1088_ _1091_ vssd1 vssd1 vccd1 vccd1 _1092_
+ sky130_fd_sc_hd__a2111o_1
X_6208_ reg_data\[16\]\[28\] _2449_ _2450_ reg_data\[9\]\[28\] vssd1 vssd1 vccd1 vccd1
+ _2778_ sky130_fd_sc_hd__a22o_1
X_7188_ reg_data\[6\]\[1\] _3131_ _3456_ vssd1 vssd1 vccd1 vccd1 _3458_ sky130_fd_sc_hd__mux2_1
X_6139_ reg_data\[20\]\[27\] _2234_ _1283_ vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__and3_1
X_9829_ clknet_leaf_50_i_clk rdata2\[13\] vssd1 vssd1 vccd1 vccd1 r_data2\[13\] sky130_fd_sc_hd__dfxtp_1
X_5510_ reg_data\[13\]\[17\] _1608_ _2102_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__and3_1
X_6490_ r_data1\[1\] _3046_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__and2_1
X_5441_ reg_data\[20\]\[16\] _1597_ _2035_ vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__and3_1
X_8160_ _3990_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__clkbuf_1
X_5372_ reg_data\[26\]\[14\] _1849_ _1850_ reg_data\[29\]\[14\] vssd1 vssd1 vccd1
+ vccd1 _1970_ sky130_fd_sc_hd__a22o_1
X_8091_ _3953_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__clkbuf_1
X_7111_ _3264_ reg_data\[8\]\[30\] _3382_ vssd1 vssd1 vccd1 vccd1 _3416_ sky130_fd_sc_hd__mux2_1
X_7042_ _3378_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__clkbuf_1
X_8993_ clknet_leaf_1_i_clk _0137_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_7944_ _3861_ reg_data\[9\]\[1\] _3859_ vssd1 vssd1 vccd1 vccd1 _3862_ sky130_fd_sc_hd__mux2_1
X_7875_ _3824_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__clkbuf_1
X_6826_ _3260_ reg_data\[22\]\[28\] _3244_ vssd1 vssd1 vccd1 vccd1 _3261_ sky130_fd_sc_hd__mux2_1
X_9614_ clknet_leaf_38_i_clk _0758_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_9545_ clknet_leaf_44_i_clk _0689_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6757_ i_data[6] vssd1 vssd1 vccd1 vccd1 _3214_ sky130_fd_sc_hd__buf_2
X_5708_ reg_data\[3\]\[20\] _1815_ _2291_ _2292_ _2293_ vssd1 vssd1 vccd1 vccd1 _2294_
+ sky130_fd_sc_hd__a2111o_1
X_6688_ _3165_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__clkbuf_1
X_9476_ clknet_leaf_63_i_clk _0620_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8427_ _4132_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__clkbuf_1
X_5639_ _2227_ vssd1 vssd1 vccd1 vccd1 rdata1\[19\] sky130_fd_sc_hd__clkbuf_1
X_8358_ _3903_ reg_data\[16\]\[21\] _4094_ vssd1 vssd1 vccd1 vccd1 _4096_ sky130_fd_sc_hd__mux2_1
X_7309_ reg_data\[5\]\[26\] _3183_ _3515_ vssd1 vssd1 vccd1 vccd1 _3522_ sky130_fd_sc_hd__mux2_1
X_8289_ _3903_ reg_data\[15\]\[21\] _4057_ vssd1 vssd1 vccd1 vccd1 _4059_ sky130_fd_sc_hd__mux2_1
X_5990_ reg_data\[1\]\[24\] _2510_ _2511_ reg_data\[15\]\[24\] vssd1 vssd1 vccd1 vccd1
+ _2568_ sky130_fd_sc_hd__a22o_1
X_4941_ reg_data\[7\]\[8\] _1081_ _1549_ _1550_ _1551_ vssd1 vssd1 vccd1 vccd1 _1552_
+ sky130_fd_sc_hd__a2111o_1
X_7660_ _3709_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__clkbuf_1
X_4872_ reg_data\[30\]\[7\] _1312_ _1313_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__and3_1
X_6611_ r_data2\[26\] _3105_ vssd1 vssd1 vccd1 vccd1 _3112_ sky130_fd_sc_hd__and2_1
X_9330_ clknet_leaf_30_i_clk _0474_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_7591_ _3672_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__clkbuf_1
X_6542_ r_data1\[26\] _3068_ vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__and2_1
X_6473_ reg_data\[7\]\[1\] _1184_ _3030_ _3031_ _3032_ vssd1 vssd1 vccd1 vccd1 _3033_
+ sky130_fd_sc_hd__a2111o_1
X_9261_ clknet_leaf_40_i_clk _0405_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_8212_ _3894_ reg_data\[14\]\[17\] _4010_ vssd1 vssd1 vccd1 vccd1 _4018_ sky130_fd_sc_hd__mux2_1
X_5424_ reg_data\[23\]\[15\] _1834_ _1835_ reg_data\[19\]\[15\] vssd1 vssd1 vccd1
+ vccd1 _2020_ sky130_fd_sc_hd__a22o_1
X_9192_ clknet_leaf_49_i_clk _0336_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_8143_ _3981_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__clkbuf_1
X_5355_ reg_data\[4\]\[14\] _1460_ _1407_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__and3_1
X_5286_ reg_data\[25\]\[13\] _1810_ _1882_ _1884_ _1885_ vssd1 vssd1 vccd1 vccd1 _1886_
+ sky130_fd_sc_hd__a2111o_1
X_8074_ _3944_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__clkbuf_1
X_7025_ reg_data\[0\]\[22\] _3175_ _3367_ vssd1 vssd1 vccd1 vccd1 _3370_ sky130_fd_sc_hd__mux2_1
X_8976_ clknet_leaf_33_i_clk _0120_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_7927_ _3851_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__clkbuf_1
X_7858_ _3814_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__clkbuf_1
X_6809_ _3249_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__clkbuf_1
X_7789_ _3256_ reg_data\[26\]\[26\] _3771_ vssd1 vssd1 vccd1 vccd1 _3778_ sky130_fd_sc_hd__mux2_1
X_9528_ clknet_leaf_13_i_clk _0672_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_9459_ clknet_leaf_30_i_clk _0603_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5140_ reg_data\[20\]\[11\] _1629_ _1743_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__and3_1
X_5071_ _1669_ _1673_ _1675_ _1677_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__or4_2
X_8830_ _4345_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__clkbuf_1
X_5973_ reg_data\[18\]\[24\] _2422_ _2120_ vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__and3_1
X_8761_ _3898_ reg_data\[29\]\[19\] _4299_ vssd1 vssd1 vccd1 vccd1 _4309_ sky130_fd_sc_hd__mux2_1
X_7712_ _3737_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__clkbuf_1
X_4924_ _1535_ vssd1 vssd1 vccd1 vccd1 rdata2\[7\] sky130_fd_sc_hd__clkbuf_1
X_8692_ _4272_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__clkbuf_1
X_4855_ reg_data\[23\]\[6\] _1206_ _1209_ reg_data\[19\]\[6\] vssd1 vssd1 vccd1 vccd1
+ _1469_ sky130_fd_sc_hd__a22o_1
X_7643_ _3246_ reg_data\[24\]\[21\] _3699_ vssd1 vssd1 vccd1 vccd1 _3701_ sky130_fd_sc_hd__mux2_1
X_4786_ _1163_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__clkbuf_4
X_7574_ reg_data\[23\]\[21\] _3173_ _3662_ vssd1 vssd1 vccd1 vccd1 _3664_ sky130_fd_sc_hd__mux2_1
X_6525_ r_data1\[18\] _3057_ vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__and2_1
X_9313_ clknet_leaf_66_i_clk _0457_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_9244_ clknet_leaf_76_i_clk _0388_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6456_ _3008_ _3012_ _3014_ _3016_ vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__or4_1
X_9175_ clknet_leaf_14_i_clk _0319_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6387_ reg_data\[5\]\[0\] _1085_ _2530_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__and3_1
X_5407_ reg_data\[25\]\[15\] _1810_ _2000_ _2001_ _2002_ vssd1 vssd1 vccd1 vccd1 _2003_
+ sky130_fd_sc_hd__a2111o_1
X_5338_ reg_data\[16\]\[14\] _1799_ _1800_ reg_data\[9\]\[14\] vssd1 vssd1 vccd1 vccd1
+ _1937_ sky130_fd_sc_hd__a22o_1
X_8126_ _3972_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__clkbuf_1
X_8057_ _3935_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__clkbuf_1
X_7008_ reg_data\[0\]\[14\] _3158_ _3356_ vssd1 vssd1 vccd1 vccd1 _3361_ sky130_fd_sc_hd__mux2_1
X_5269_ reg_data\[14\]\[13\] _1608_ _1090_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__and3_1
X_8959_ clknet_leaf_73_i_clk _0103_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_4640_ reg_data\[23\]\[3\] _1099_ _1101_ reg_data\[19\]\[3\] vssd1 vssd1 vccd1 vccd1
+ _1261_ sky130_fd_sc_hd__a22o_1
X_6310_ reg_data\[7\]\[30\] _2433_ _2873_ _2874_ _2875_ vssd1 vssd1 vccd1 vccd1 _2876_
+ sky130_fd_sc_hd__a2111o_1
X_4571_ _1163_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__buf_2
X_7290_ reg_data\[5\]\[17\] _3164_ _3504_ vssd1 vssd1 vccd1 vccd1 _3512_ sky130_fd_sc_hd__mux2_1
X_6241_ reg_data\[22\]\[29\] _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__and3_1
X_6172_ reg_data\[14\]\[28\] _2473_ _2156_ vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__and3_1
X_5123_ reg_data\[2\]\[11\] _1613_ _1104_ _1106_ reg_data\[11\]\[11\] vssd1 vssd1
+ vccd1 vccd1 _1728_ sky130_fd_sc_hd__a32o_1
X_5054_ reg_data\[6\]\[10\] _1600_ _1048_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__and3_1
X_9862_ clknet_leaf_72_i_clk _0932_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_8813_ reg_data\[11\]\[11\] i_data[11] _4335_ vssd1 vssd1 vccd1 vccd1 _4337_ sky130_fd_sc_hd__mux2_1
X_9793_ clknet_leaf_72_i_clk rdata1\[9\] vssd1 vssd1 vccd1 vccd1 r_data1\[9\] sky130_fd_sc_hd__dfxtp_1
X_5956_ reg_data\[13\]\[24\] _2214_ _2102_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__and3_1
X_8744_ _4300_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__clkbuf_1
X_5887_ reg_data\[6\]\[23\] _2207_ _2323_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__and3_1
X_8675_ reg_data\[19\]\[10\] _3149_ _4263_ vssd1 vssd1 vccd1 vccd1 _4264_ sky130_fd_sc_hd__mux2_1
X_4907_ reg_data\[4\]\[7\] _1460_ _1407_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__and3_1
X_7626_ _3229_ reg_data\[24\]\[13\] _3688_ vssd1 vssd1 vccd1 vccd1 _3692_ sky130_fd_sc_hd__mux2_1
X_4838_ reg_data\[21\]\[6\] _1272_ _1273_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__and3_1
X_7557_ reg_data\[23\]\[13\] _3156_ _3651_ vssd1 vssd1 vccd1 vccd1 _3655_ sky130_fd_sc_hd__mux2_1
X_4769_ reg_data\[23\]\[5\] _1099_ _1101_ reg_data\[19\]\[5\] vssd1 vssd1 vccd1 vccd1
+ _1386_ sky130_fd_sc_hd__a22o_1
X_6508_ _3045_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__clkbuf_2
X_7488_ _3229_ reg_data\[21\]\[13\] _3614_ vssd1 vssd1 vccd1 vccd1 _3618_ sky130_fd_sc_hd__mux2_1
X_6439_ reg_data\[6\]\[1\] _1020_ _1236_ vssd1 vssd1 vccd1 vccd1 _3000_ sky130_fd_sc_hd__and3_1
X_9227_ clknet_leaf_44_i_clk _0371_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_9158_ clknet_leaf_47_i_clk _0302_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8109_ _3857_ reg_data\[13\]\[0\] _3963_ vssd1 vssd1 vccd1 vccd1 _3964_ sky130_fd_sc_hd__mux2_1
X_9089_ clknet_leaf_2_i_clk _0233_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_50_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5810_ _1098_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__buf_2
X_6790_ _3236_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__clkbuf_1
X_5741_ reg_data\[4\]\[21\] _2325_ _1863_ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__and3_1
X_8460_ _3869_ reg_data\[18\]\[5\] _4144_ vssd1 vssd1 vccd1 vccd1 _4150_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_65_i_clk clknet_3_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5672_ reg_data\[21\]\[20\] _2086_ _2087_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__and3_1
X_7411_ _3564_ vssd1 vssd1 vccd1 vccd1 _3576_ sky130_fd_sc_hd__buf_4
X_4623_ reg_data\[20\]\[3\] _1058_ _1060_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__and3_1
X_8391_ _4113_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__clkbuf_1
X_4554_ reg_data\[5\]\[2\] _1175_ _1144_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__and3_1
X_7342_ _3539_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__clkbuf_1
X_7273_ reg_data\[5\]\[9\] _3147_ _3493_ vssd1 vssd1 vccd1 vccd1 _3503_ sky130_fd_sc_hd__mux2_1
X_9012_ clknet_leaf_18_i_clk _0156_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6224_ reg_data\[5\]\[29\] _1085_ _2530_ vssd1 vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__and3_1
X_4485_ _1040_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__buf_4
X_6155_ reg_data\[8\]\[27\] _2447_ _2448_ reg_data\[10\]\[27\] _2726_ vssd1 vssd1
+ vccd1 vccd1 _2727_ sky130_fd_sc_hd__a221o_1
X_6086_ reg_data\[3\]\[26\] _2421_ _2657_ _2658_ _2659_ vssd1 vssd1 vccd1 vccd1 _2660_
+ sky130_fd_sc_hd__a2111o_1
X_5106_ reg_data\[25\]\[11\] _1037_ _1707_ _1709_ _1710_ vssd1 vssd1 vccd1 vccd1 _1711_
+ sky130_fd_sc_hd__a2111o_1
X_9914_ clknet_leaf_32_i_clk _0984_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_5037_ reg_data\[27\]\[9\] _1199_ _1642_ _1643_ _1644_ vssd1 vssd1 vccd1 vccd1 _1645_
+ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_18_i_clk clknet_3_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_9845_ clknet_leaf_39_i_clk rdata2\[29\] vssd1 vssd1 vccd1 vccd1 r_data2\[29\] sky130_fd_sc_hd__dfxtp_1
X_9776_ clknet_leaf_35_i_clk _0920_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_8727_ _4291_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__clkbuf_1
X_6988_ _3350_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__clkbuf_1
X_5939_ _2518_ vssd1 vssd1 vccd1 vccd1 rdata2\[23\] sky130_fd_sc_hd__clkbuf_1
X_8658_ reg_data\[19\]\[2\] _3133_ _4252_ vssd1 vssd1 vccd1 vccd1 _4255_ sky130_fd_sc_hd__mux2_1
X_8589_ _4218_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__clkbuf_1
X_7609_ _3212_ reg_data\[24\]\[5\] _3677_ vssd1 vssd1 vccd1 vccd1 _3683_ sky130_fd_sc_hd__mux2_1
X_7960_ _3872_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__clkbuf_1
X_6911_ _3195_ reg_data\[10\]\[0\] _3309_ vssd1 vssd1 vccd1 vccd1 _3310_ sky130_fd_sc_hd__mux2_1
X_7891_ _3832_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__clkbuf_1
X_6842_ _3272_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__clkbuf_1
X_9630_ clknet_leaf_7_i_clk _0774_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6773_ i_data[11] vssd1 vssd1 vccd1 vccd1 _3225_ sky130_fd_sc_hd__buf_2
X_9561_ clknet_leaf_72_i_clk _0705_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_9492_ clknet_leaf_18_i_clk _0636_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_8512_ _3921_ reg_data\[18\]\[30\] _4143_ vssd1 vssd1 vccd1 vccd1 _4177_ sky130_fd_sc_hd__mux2_1
X_5724_ reg_data\[16\]\[20\] _1843_ _1844_ reg_data\[9\]\[20\] vssd1 vssd1 vccd1 vccd1
+ _2310_ sky130_fd_sc_hd__a22o_1
X_8443_ _4140_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__clkbuf_1
X_5655_ reg_data\[12\]\[19\] _1693_ _1187_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__and3_1
X_8374_ _3919_ reg_data\[16\]\[29\] _4094_ vssd1 vssd1 vccd1 vccd1 _4104_ sky130_fd_sc_hd__mux2_1
X_4606_ _1227_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__clkbuf_4
X_5586_ reg_data\[20\]\[18\] _2005_ _1342_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__and3_1
X_7325_ reg_data\[3\]\[1\] _3131_ _3529_ vssd1 vssd1 vccd1 vccd1 _3531_ sky130_fd_sc_hd__mux2_1
X_4537_ _1142_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__buf_2
X_7256_ _3494_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__clkbuf_1
X_4468_ reg_data\[14\]\[2\] _1089_ _1090_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__and3_1
X_6207_ reg_data\[27\]\[28\] _2439_ _2774_ _2775_ _2776_ vssd1 vssd1 vccd1 vccd1 _2777_
+ sky130_fd_sc_hd__a2111o_1
X_7187_ _3457_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__clkbuf_1
X_6138_ reg_data\[30\]\[27\] _1146_ _2006_ vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__and3_1
X_4399_ _0994_ rs1\[1\] _1023_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__a2bb2o_1
X_6069_ reg_data\[23\]\[26\] _2393_ _2394_ reg_data\[19\]\[26\] vssd1 vssd1 vccd1
+ vccd1 _2644_ sky130_fd_sc_hd__a22o_1
X_9828_ clknet_leaf_50_i_clk rdata2\[12\] vssd1 vssd1 vccd1 vccd1 r_data2\[12\] sky130_fd_sc_hd__dfxtp_1
X_9759_ clknet_leaf_0_i_clk _0903_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5440_ _1059_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__clkbuf_4
X_5371_ reg_data\[8\]\[14\] _1841_ _1842_ reg_data\[10\]\[14\] _1968_ vssd1 vssd1
+ vccd1 vccd1 _1969_ sky130_fd_sc_hd__a221o_1
X_8090_ _3909_ reg_data\[30\]\[24\] _3948_ vssd1 vssd1 vccd1 vccd1 _3953_ sky130_fd_sc_hd__mux2_1
X_7110_ _3415_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
X_7041_ reg_data\[0\]\[30\] _3191_ _3344_ vssd1 vssd1 vccd1 vccd1 _3378_ sky130_fd_sc_hd__mux2_1
X_8992_ clknet_leaf_1_i_clk _0136_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7943_ i_data[1] vssd1 vssd1 vccd1 vccd1 _3861_ sky130_fd_sc_hd__clkbuf_4
X_7874_ _3204_ reg_data\[28\]\[1\] _3822_ vssd1 vssd1 vccd1 vccd1 _3824_ sky130_fd_sc_hd__mux2_1
X_6825_ i_data[28] vssd1 vssd1 vccd1 vccd1 _3260_ sky130_fd_sc_hd__clkbuf_4
X_9613_ clknet_leaf_50_i_clk _0757_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6756_ _3213_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__clkbuf_1
X_9544_ clknet_leaf_46_i_clk _0688_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_5707_ reg_data\[30\]\[20\] _2234_ _1344_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__and3_1
X_6687_ reg_data\[4\]\[17\] _3164_ _3150_ vssd1 vssd1 vccd1 vccd1 _3165_ sky130_fd_sc_hd__mux2_1
X_9475_ clknet_leaf_65_i_clk _0619_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8426_ _3903_ reg_data\[17\]\[21\] _4130_ vssd1 vssd1 vccd1 vccd1 _4132_ sky130_fd_sc_hd__mux2_1
X_5638_ _2217_ _2222_ _2224_ _2226_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__or4_1
X_5569_ reg_data\[7\]\[18\] _1780_ _2157_ _2158_ _2159_ vssd1 vssd1 vccd1 vccd1 _2160_
+ sky130_fd_sc_hd__a2111o_1
X_8357_ _4095_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__clkbuf_1
X_7308_ _3521_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__clkbuf_1
X_8288_ _4058_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__clkbuf_1
X_7239_ _3484_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__clkbuf_1
X_4940_ reg_data\[13\]\[8\] _1089_ _1257_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__and3_1
X_4871_ reg_data\[18\]\[7\] _1055_ _1483_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__and3_1
X_7590_ reg_data\[23\]\[29\] _3189_ _3662_ vssd1 vssd1 vccd1 vccd1 _3672_ sky130_fd_sc_hd__mux2_1
X_6610_ _3111_ vssd1 vssd1 vccd1 vccd1 o_data2[25] sky130_fd_sc_hd__buf_2
X_6541_ _3074_ vssd1 vssd1 vccd1 vccd1 o_data1[25] sky130_fd_sc_hd__buf_2
X_6472_ reg_data\[12\]\[1\] _2562_ _1289_ vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__and3_1
X_9260_ clknet_leaf_40_i_clk _0404_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_9191_ clknet_leaf_48_i_clk _0335_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_5423_ _2003_ _2009_ _2013_ _2018_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__or4_1
X_8211_ _4017_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__clkbuf_1
X_5354_ reg_data\[6\]\[14\] _1951_ _1632_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__and3_1
X_8142_ _3892_ reg_data\[13\]\[16\] _3974_ vssd1 vssd1 vccd1 vccd1 _3981_ sky130_fd_sc_hd__mux2_1
X_5285_ reg_data\[22\]\[13\] _1509_ _1152_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__and3_1
X_8073_ _3892_ reg_data\[30\]\[16\] _3937_ vssd1 vssd1 vccd1 vccd1 _3944_ sky130_fd_sc_hd__mux2_1
X_7024_ _3369_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__clkbuf_1
X_8975_ clknet_leaf_32_i_clk _0119_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_7926_ _3256_ reg_data\[28\]\[26\] _3844_ vssd1 vssd1 vccd1 vccd1 _3851_ sky130_fd_sc_hd__mux2_1
X_7857_ _3256_ reg_data\[27\]\[26\] _3807_ vssd1 vssd1 vccd1 vccd1 _3814_ sky130_fd_sc_hd__mux2_1
X_6808_ _3248_ reg_data\[22\]\[22\] _3244_ vssd1 vssd1 vccd1 vccd1 _3249_ sky130_fd_sc_hd__mux2_1
X_7788_ _3777_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__clkbuf_1
X_9527_ clknet_leaf_13_i_clk _0671_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6739_ _3201_ vssd1 vssd1 vccd1 vccd1 _3202_ sky130_fd_sc_hd__buf_4
X_9458_ clknet_leaf_31_i_clk _0602_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_8409_ _3886_ reg_data\[17\]\[13\] _4119_ vssd1 vssd1 vccd1 vccd1 _4123_ sky130_fd_sc_hd__mux2_1
X_9389_ clknet_leaf_40_i_clk _0533_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5070_ reg_data\[24\]\[10\] _1127_ _1130_ reg_data\[28\]\[10\] _1676_ vssd1 vssd1
+ vccd1 vccd1 _1677_ sky130_fd_sc_hd__a221o_1
X_5972_ reg_data\[25\]\[24\] _2416_ _2547_ _2548_ _2549_ vssd1 vssd1 vccd1 vccd1 _2550_
+ sky130_fd_sc_hd__a2111o_1
X_8760_ _4308_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__clkbuf_1
X_7711_ _3246_ reg_data\[25\]\[21\] _3735_ vssd1 vssd1 vccd1 vccd1 _3737_ sky130_fd_sc_hd__mux2_1
X_4923_ _1526_ _1530_ _1532_ _1534_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__or4_1
X_8691_ reg_data\[19\]\[18\] _3166_ _4263_ vssd1 vssd1 vccd1 vccd1 _4272_ sky130_fd_sc_hd__mux2_1
X_4854_ _1454_ _1458_ _1463_ _1467_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__or4_1
X_7642_ _3700_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__clkbuf_1
X_4785_ _1138_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__buf_2
X_7573_ _3663_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__clkbuf_1
X_6524_ _3065_ vssd1 vssd1 vccd1 vccd1 o_data1[17] sky130_fd_sc_hd__buf_2
X_9312_ clknet_leaf_66_i_clk _0456_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_9243_ clknet_leaf_76_i_clk _0387_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6455_ reg_data\[24\]\[1\] _1126_ _1129_ reg_data\[28\]\[1\] _3015_ vssd1 vssd1 vccd1
+ vccd1 _3016_ sky130_fd_sc_hd__a221o_1
X_9174_ clknet_leaf_15_i_clk _0318_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6386_ reg_data\[4\]\[0\] _1072_ _2469_ vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__and3_1
X_5406_ reg_data\[21\]\[15\] _1509_ _1510_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__and3_1
X_5337_ reg_data\[27\]\[14\] _1786_ _1933_ _1934_ _1935_ vssd1 vssd1 vccd1 vccd1 _1936_
+ sky130_fd_sc_hd__a2111o_1
X_8125_ _3875_ reg_data\[13\]\[8\] _3963_ vssd1 vssd1 vccd1 vccd1 _3972_ sky130_fd_sc_hd__mux2_1
X_8056_ _3875_ reg_data\[30\]\[8\] _3926_ vssd1 vssd1 vccd1 vccd1 _3935_ sky130_fd_sc_hd__mux2_1
X_5268_ reg_data\[12\]\[13\] _1381_ _1606_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__and3_1
X_7007_ _3360_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__clkbuf_1
X_5199_ reg_data\[8\]\[12\] _1797_ _1798_ reg_data\[10\]\[12\] _1801_ vssd1 vssd1
+ vccd1 vccd1 _1802_ sky130_fd_sc_hd__a221o_1
X_8958_ clknet_leaf_74_i_clk _0102_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_7909_ _3239_ reg_data\[28\]\[18\] _3833_ vssd1 vssd1 vccd1 vccd1 _3842_ sky130_fd_sc_hd__mux2_1
X_8889_ clknet_leaf_9_i_clk _0033_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_4570_ reg_data\[13\]\[2\] _1189_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__and3_1
X_6240_ _2808_ vssd1 vssd1 vccd1 vccd1 rdata1\[29\] sky130_fd_sc_hd__clkbuf_1
X_6171_ reg_data\[0\]\[28\] _2381_ _2739_ _2740_ _2741_ vssd1 vssd1 vccd1 vccd1 _2742_
+ sky130_fd_sc_hd__a2111o_1
X_5122_ reg_data\[23\]\[11\] _1099_ _1101_ reg_data\[19\]\[11\] vssd1 vssd1 vccd1
+ vccd1 _1727_ sky130_fd_sc_hd__a22o_1
X_5053_ reg_data\[3\]\[10\] _1054_ _1657_ _1658_ _1659_ vssd1 vssd1 vccd1 vccd1 _1660_
+ sky130_fd_sc_hd__a2111o_1
X_9861_ clknet_leaf_71_i_clk _0931_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_8812_ _4336_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__clkbuf_1
X_9792_ clknet_leaf_55_i_clk rdata1\[8\] vssd1 vssd1 vccd1 vccd1 r_data1\[8\] sky130_fd_sc_hd__dfxtp_1
X_5955_ reg_data\[12\]\[24\] _1986_ _2271_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__and3_1
X_8743_ _3879_ reg_data\[29\]\[10\] _4299_ vssd1 vssd1 vccd1 vccd1 _4300_ sky130_fd_sc_hd__mux2_1
X_5886_ reg_data\[3\]\[23\] _2376_ _2464_ _2465_ _2466_ vssd1 vssd1 vccd1 vccd1 _2467_
+ sky130_fd_sc_hd__a2111o_1
X_8674_ _4251_ vssd1 vssd1 vccd1 vccd1 _4263_ sky130_fd_sc_hd__buf_4
X_4906_ reg_data\[6\]\[7\] _1347_ _1152_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__and3_1
X_7625_ _3691_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__clkbuf_1
X_4837_ reg_data\[22\]\[6\] _1143_ _1270_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__and3_1
X_7556_ _3654_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__clkbuf_1
X_4768_ _1370_ _1374_ _1378_ _1384_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__or4_2
X_6507_ _3056_ vssd1 vssd1 vccd1 vccd1 o_data1[9] sky130_fd_sc_hd__buf_2
X_7487_ _3617_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__clkbuf_1
X_4699_ reg_data\[6\]\[4\] _1072_ _1048_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__and3_1
X_9226_ clknet_leaf_41_i_clk _0370_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6438_ reg_data\[3\]\[1\] _1053_ _2996_ _2997_ _2998_ vssd1 vssd1 vccd1 vccd1 _2999_
+ sky130_fd_sc_hd__a2111o_1
X_9157_ clknet_leaf_62_i_clk _0301_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6369_ reg_data\[1\]\[31\] _2510_ _2511_ reg_data\[15\]\[31\] vssd1 vssd1 vccd1 vccd1
+ _2933_ sky130_fd_sc_hd__a22o_1
X_8108_ _3962_ vssd1 vssd1 vccd1 vccd1 _3963_ sky130_fd_sc_hd__buf_4
X_9088_ clknet_leaf_0_i_clk _0232_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8039_ _3925_ vssd1 vssd1 vccd1 vccd1 _3926_ sky130_fd_sc_hd__buf_4
X_5740_ _1071_ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__buf_2
X_5671_ reg_data\[17\]\[20\] _1766_ _1708_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__and3_1
X_7410_ _3575_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__clkbuf_1
X_4622_ reg_data\[18\]\[3\] _1055_ _1064_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__and3_1
X_8390_ _3867_ reg_data\[17\]\[4\] _4108_ vssd1 vssd1 vccd1 vccd1 _4113_ sky130_fd_sc_hd__mux2_1
X_4553_ _0999_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__clkbuf_4
X_7341_ reg_data\[3\]\[9\] _3147_ _3529_ vssd1 vssd1 vccd1 vccd1 _3539_ sky130_fd_sc_hd__mux2_1
X_4484_ reg_data\[2\]\[2\] _1103_ _1104_ _1106_ reg_data\[11\]\[2\] vssd1 vssd1 vccd1
+ vccd1 _1107_ sky130_fd_sc_hd__a32o_1
X_7272_ _3502_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__clkbuf_1
X_9011_ clknet_leaf_18_i_clk _0155_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6223_ reg_data\[4\]\[29\] _2325_ _2469_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__and3_1
X_6154_ reg_data\[16\]\[27\] _2449_ _2450_ reg_data\[9\]\[27\] vssd1 vssd1 vccd1 vccd1
+ _2726_ sky130_fd_sc_hd__a22o_1
X_6085_ reg_data\[20\]\[26\] _2234_ _1283_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__and3_1
X_5105_ reg_data\[21\]\[11\] _1480_ _1240_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__and3_1
X_9913_ clknet_leaf_37_i_clk _0983_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_5036_ reg_data\[1\]\[9\] _1298_ _1299_ reg_data\[15\]\[9\] vssd1 vssd1 vccd1 vccd1
+ _1644_ sky130_fd_sc_hd__a22o_1
X_9844_ clknet_leaf_32_i_clk rdata2\[28\] vssd1 vssd1 vccd1 vccd1 r_data2\[28\] sky130_fd_sc_hd__dfxtp_1
X_9775_ clknet_leaf_37_i_clk _0919_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6987_ reg_data\[0\]\[4\] _3137_ _3345_ vssd1 vssd1 vccd1 vccd1 _3350_ sky130_fd_sc_hd__mux2_1
X_5938_ _2505_ _2513_ _2515_ _2517_ vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__or4_1
X_8726_ _3863_ reg_data\[29\]\[2\] _4288_ vssd1 vssd1 vccd1 vccd1 _4291_ sky130_fd_sc_hd__mux2_1
X_5869_ reg_data\[16\]\[22\] _2449_ _2450_ reg_data\[9\]\[22\] vssd1 vssd1 vccd1 vccd1
+ _2451_ sky130_fd_sc_hd__a22o_1
X_8657_ _4254_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__clkbuf_1
X_8588_ _3861_ reg_data\[12\]\[1\] _4216_ vssd1 vssd1 vccd1 vccd1 _4218_ sky130_fd_sc_hd__mux2_1
X_7608_ _3682_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__clkbuf_1
X_7539_ _3645_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__clkbuf_1
X_9209_ clknet_leaf_8_i_clk _0353_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_7890_ _3220_ reg_data\[28\]\[9\] _3822_ vssd1 vssd1 vccd1 vccd1 _3832_ sky130_fd_sc_hd__mux2_1
X_6910_ _3308_ vssd1 vssd1 vccd1 vccd1 _3309_ sky130_fd_sc_hd__buf_4
X_6841_ reg_data\[2\]\[0\] _3118_ _3271_ vssd1 vssd1 vccd1 vccd1 _3272_ sky130_fd_sc_hd__mux2_1
X_9560_ clknet_leaf_68_i_clk _0704_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8511_ _4176_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__clkbuf_1
X_6772_ _3224_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__clkbuf_1
X_9491_ clknet_leaf_18_i_clk _0635_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5723_ reg_data\[27\]\[20\] _1833_ _2306_ _2307_ _2308_ vssd1 vssd1 vccd1 vccd1 _2309_
+ sky130_fd_sc_hd__a2111o_1
X_8442_ _3919_ reg_data\[17\]\[29\] _4130_ vssd1 vssd1 vccd1 vccd1 _4140_ sky130_fd_sc_hd__mux2_1
X_5654_ reg_data\[14\]\[19\] _2183_ _1164_ vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__and3_1
X_8373_ _4103_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__clkbuf_1
X_4605_ _1166_ _1226_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__and2_2
X_5585_ reg_data\[18\]\[18\] _1816_ _2120_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__and3_1
X_7324_ _3530_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__clkbuf_1
X_4536_ _1157_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__clkbuf_4
X_4467_ _1056_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__clkbuf_4
X_7255_ reg_data\[5\]\[0\] _3118_ _3493_ vssd1 vssd1 vccd1 vccd1 _3494_ sky130_fd_sc_hd__mux2_1
X_6206_ reg_data\[1\]\[28\] _2510_ _2511_ reg_data\[15\]\[28\] vssd1 vssd1 vccd1 vccd1
+ _2776_ sky130_fd_sc_hd__a22o_1
X_4398_ i_rs1[0] i_rs1[1] i_rs_valid vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__o21a_1
X_7186_ reg_data\[6\]\[0\] _3118_ _3456_ vssd1 vssd1 vccd1 vccd1 _3457_ sky130_fd_sc_hd__mux2_1
X_6137_ reg_data\[18\]\[27\] _2422_ _1167_ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__and3_1
X_6068_ _2630_ _2634_ _2638_ _2642_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__or4_2
X_5019_ reg_data\[18\]\[9\] _1159_ _1513_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__and3_1
X_9827_ clknet_leaf_59_i_clk rdata2\[11\] vssd1 vssd1 vccd1 vccd1 r_data2\[11\] sky130_fd_sc_hd__dfxtp_1
X_9758_ clknet_leaf_77_i_clk _0902_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8709_ _4281_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__clkbuf_1
X_9689_ clknet_leaf_72_i_clk _0833_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_64_i_clk clknet_3_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_17_i_clk clknet_3_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5370_ reg_data\[16\]\[14\] _1843_ _1844_ reg_data\[9\]\[14\] vssd1 vssd1 vccd1 vccd1
+ _1968_ sky130_fd_sc_hd__a22o_1
X_7040_ _3377_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__clkbuf_1
X_8991_ clknet_leaf_2_i_clk _0135_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_7942_ _3860_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__clkbuf_1
X_7873_ _3823_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__clkbuf_1
X_9612_ clknet_leaf_50_i_clk _0756_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6824_ _3259_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__clkbuf_1
X_6755_ _3212_ reg_data\[22\]\[5\] _3202_ vssd1 vssd1 vccd1 vccd1 _3213_ sky130_fd_sc_hd__mux2_1
X_9543_ clknet_leaf_26_i_clk _0687_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_5706_ reg_data\[20\]\[20\] _2005_ _1342_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__and3_1
X_9474_ clknet_leaf_66_i_clk _0618_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8425_ _4131_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__clkbuf_1
X_6686_ i_data[17] vssd1 vssd1 vccd1 vccd1 _3164_ sky130_fd_sc_hd__clkbuf_4
X_5637_ reg_data\[24\]\[19\] _1803_ _1804_ reg_data\[28\]\[19\] _2225_ vssd1 vssd1
+ vccd1 vccd1 _2226_ sky130_fd_sc_hd__a221o_1
X_5568_ reg_data\[13\]\[18\] _1608_ _2102_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__and3_1
X_8356_ _3900_ reg_data\[16\]\[20\] _4094_ vssd1 vssd1 vccd1 vccd1 _4095_ sky130_fd_sc_hd__mux2_1
X_7307_ reg_data\[5\]\[25\] _3181_ _3515_ vssd1 vssd1 vccd1 vccd1 _3521_ sky130_fd_sc_hd__mux2_1
X_8287_ _3900_ reg_data\[15\]\[20\] _4057_ vssd1 vssd1 vccd1 vccd1 _4058_ sky130_fd_sc_hd__mux2_1
X_4519_ _1140_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__clkbuf_4
X_7238_ reg_data\[6\]\[25\] _3181_ _3478_ vssd1 vssd1 vccd1 vccd1 _3484_ sky130_fd_sc_hd__mux2_1
X_5499_ reg_data\[30\]\[17\] _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__and3_1
X_7169_ _3447_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__clkbuf_1
X_4870_ _1063_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__clkbuf_4
X_6540_ r_data1\[25\] _3068_ vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__and2_1
X_6471_ reg_data\[14\]\[1\] _1186_ _1344_ vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__and3_1
X_9190_ clknet_leaf_48_i_clk _0334_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_5422_ reg_data\[7\]\[15\] _1827_ _2014_ _2015_ _2017_ vssd1 vssd1 vccd1 vccd1 _2018_
+ sky130_fd_sc_hd__a2111o_1
X_8210_ _3892_ reg_data\[14\]\[16\] _4010_ vssd1 vssd1 vccd1 vccd1 _4017_ sky130_fd_sc_hd__mux2_1
X_5353_ _0999_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__clkbuf_4
X_8141_ _3980_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__clkbuf_1
X_5284_ reg_data\[21\]\[13\] _1883_ _1273_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__and3_1
X_8072_ _3943_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__clkbuf_1
X_7023_ reg_data\[0\]\[21\] _3173_ _3367_ vssd1 vssd1 vccd1 vccd1 _3369_ sky130_fd_sc_hd__mux2_1
X_8974_ clknet_leaf_37_i_clk _0118_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_7925_ _3850_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__clkbuf_1
X_7856_ _3813_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__clkbuf_1
X_6807_ i_data[22] vssd1 vssd1 vccd1 vccd1 _3248_ sky130_fd_sc_hd__buf_2
X_7787_ _3254_ reg_data\[26\]\[25\] _3771_ vssd1 vssd1 vccd1 vccd1 _3777_ sky130_fd_sc_hd__mux2_1
X_9526_ clknet_leaf_14_i_clk _0670_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_4999_ _1067_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__buf_2
X_6738_ _3198_ _3200_ vssd1 vssd1 vccd1 vccd1 _3201_ sky130_fd_sc_hd__nand2_2
X_9457_ clknet_leaf_31_i_clk _0601_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6669_ reg_data\[4\]\[11\] _3152_ _3150_ vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__mux2_1
X_9388_ clknet_leaf_39_i_clk _0532_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8408_ _4122_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__clkbuf_1
X_8339_ _3884_ reg_data\[16\]\[12\] _4083_ vssd1 vssd1 vccd1 vccd1 _4086_ sky130_fd_sc_hd__mux2_1
X_5971_ reg_data\[17\]\[24\] _2117_ _1148_ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__and3_1
X_7710_ _3736_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__clkbuf_1
X_8690_ _4271_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__clkbuf_1
X_4922_ reg_data\[24\]\[7\] _1225_ _1228_ reg_data\[28\]\[7\] _1533_ vssd1 vssd1 vccd1
+ vccd1 _1534_ sky130_fd_sc_hd__a221o_1
X_7641_ _3243_ reg_data\[24\]\[20\] _3699_ vssd1 vssd1 vccd1 vccd1 _3700_ sky130_fd_sc_hd__mux2_1
X_4853_ reg_data\[7\]\[6\] _1185_ _1464_ _1465_ _1466_ vssd1 vssd1 vccd1 vccd1 _1467_
+ sky130_fd_sc_hd__a2111o_1
X_4784_ reg_data\[18\]\[5\] _1159_ _1168_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__and3_1
X_7572_ reg_data\[23\]\[20\] _3170_ _3662_ vssd1 vssd1 vccd1 vccd1 _3663_ sky130_fd_sc_hd__mux2_1
X_6523_ r_data1\[17\] _3057_ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__and2_1
X_9311_ clknet_leaf_67_i_clk _0455_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_9242_ clknet_leaf_74_i_clk _0386_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6454_ reg_data\[26\]\[1\] _1131_ _1133_ reg_data\[29\]\[1\] vssd1 vssd1 vccd1 vccd1
+ _3015_ sky130_fd_sc_hd__a22o_1
X_5405_ reg_data\[17\]\[15\] _1883_ _1395_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__and3_1
X_9173_ clknet_leaf_20_i_clk _0317_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6385_ reg_data\[6\]\[0\] _1020_ _1236_ vssd1 vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__and3_1
X_5336_ reg_data\[1\]\[14\] _1729_ _1793_ _1794_ reg_data\[15\]\[14\] vssd1 vssd1
+ vccd1 vccd1 _1935_ sky130_fd_sc_hd__a32o_1
X_8124_ _3971_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__clkbuf_1
X_8055_ _3934_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__clkbuf_1
X_5267_ reg_data\[13\]\[13\] _1867_ _1087_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__and3_1
X_7006_ reg_data\[0\]\[13\] _3156_ _3356_ vssd1 vssd1 vccd1 vccd1 _3360_ sky130_fd_sc_hd__mux2_1
X_5198_ reg_data\[16\]\[12\] _1799_ _1800_ reg_data\[9\]\[12\] vssd1 vssd1 vccd1 vccd1
+ _1801_ sky130_fd_sc_hd__a22o_1
X_8957_ clknet_leaf_71_i_clk _0101_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_7908_ _3841_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__clkbuf_1
X_8888_ clknet_leaf_9_i_clk _0032_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_7839_ _3804_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__clkbuf_1
X_9509_ clknet_leaf_65_i_clk _0653_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6170_ reg_data\[5\]\[28\] _1085_ _2530_ vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__and3_1
X_5121_ _1711_ _1715_ _1721_ _1725_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__or4_1
X_5052_ reg_data\[20\]\[10\] _1597_ _1315_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__and3_1
X_9860_ clknet_leaf_70_i_clk _0930_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_9791_ clknet_leaf_55_i_clk rdata1\[7\] vssd1 vssd1 vccd1 vccd1 r_data1\[7\] sky130_fd_sc_hd__dfxtp_1
X_8811_ reg_data\[11\]\[10\] i_data[10] _4335_ vssd1 vssd1 vccd1 vccd1 _4336_ sky130_fd_sc_hd__mux2_1
X_8742_ _4287_ vssd1 vssd1 vccd1 vccd1 _4299_ sky130_fd_sc_hd__buf_4
X_5954_ reg_data\[14\]\[24\] _2473_ _2156_ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__and3_1
X_5885_ reg_data\[20\]\[23\] _2204_ _2035_ vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__and3_1
X_8673_ _4262_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__clkbuf_1
X_4905_ reg_data\[3\]\[7\] _1158_ _1514_ _1515_ _1516_ vssd1 vssd1 vccd1 vccd1 _1517_
+ sky130_fd_sc_hd__a2111o_1
X_4836_ _1450_ vssd1 vssd1 vccd1 vccd1 rdata1\[6\] sky130_fd_sc_hd__clkbuf_2
X_7624_ _3227_ reg_data\[24\]\[12\] _3688_ vssd1 vssd1 vccd1 vccd1 _3691_ sky130_fd_sc_hd__mux2_1
X_7555_ reg_data\[23\]\[12\] _3154_ _3651_ vssd1 vssd1 vccd1 vccd1 _3654_ sky130_fd_sc_hd__mux2_1
X_6506_ r_data1\[9\] _3046_ vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__and2_1
X_4767_ reg_data\[7\]\[5\] _1081_ _1380_ _1382_ _1383_ vssd1 vssd1 vccd1 vccd1 _1384_
+ sky130_fd_sc_hd__a2111o_1
X_7486_ _3227_ reg_data\[21\]\[12\] _3614_ vssd1 vssd1 vccd1 vccd1 _3617_ sky130_fd_sc_hd__mux2_1
X_4698_ reg_data\[3\]\[4\] _1054_ _1311_ _1314_ _1316_ vssd1 vssd1 vccd1 vccd1 _1317_
+ sky130_fd_sc_hd__a2111o_1
X_6437_ reg_data\[20\]\[1\] _1046_ _1248_ vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__and3_1
X_9225_ clknet_leaf_49_i_clk _0369_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6368_ reg_data\[2\]\[31\] _2443_ _2507_ _2508_ reg_data\[11\]\[31\] vssd1 vssd1
+ vccd1 vccd1 _2932_ sky130_fd_sc_hd__a32o_1
X_9156_ clknet_leaf_63_i_clk _0300_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_5319_ _1034_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__buf_2
X_8107_ _3601_ _3961_ vssd1 vssd1 vccd1 vccd1 _3962_ sky130_fd_sc_hd__nand2_2
X_6299_ reg_data\[18\]\[30\] _2422_ _1167_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__and3_1
X_9087_ clknet_leaf_0_i_clk _0231_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8038_ _3268_ _3820_ vssd1 vssd1 vccd1 vccd1 _3925_ sky130_fd_sc_hd__or2_2
X_5670_ reg_data\[22\]\[20\] _2143_ _2256_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__and3_1
X_4621_ reg_data\[25\]\[3\] _1037_ _1237_ _1239_ _1241_ vssd1 vssd1 vccd1 vccd1 _1242_
+ sky130_fd_sc_hd__a2111o_1
X_4552_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__buf_4
X_7340_ _3538_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__clkbuf_1
X_4483_ _1105_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__buf_4
X_7271_ reg_data\[5\]\[8\] _3145_ _3493_ vssd1 vssd1 vccd1 vccd1 _3502_ sky130_fd_sc_hd__mux2_1
X_9010_ clknet_leaf_17_i_clk _0154_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6222_ reg_data\[6\]\[29\] _1020_ _2323_ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__and3_1
X_6153_ reg_data\[27\]\[27\] _2439_ _2722_ _2723_ _2724_ vssd1 vssd1 vccd1 vccd1 _2725_
+ sky130_fd_sc_hd__a2111o_1
X_6084_ reg_data\[30\]\[26\] _1146_ _2006_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__and3_1
X_5104_ reg_data\[17\]\[11\] _1042_ _1708_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__and3_1
X_9912_ clknet_leaf_39_i_clk _0982_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_5035_ reg_data\[2\]\[9\] _1002_ _1295_ _1296_ reg_data\[11\]\[9\] vssd1 vssd1 vccd1
+ vccd1 _1643_ sky130_fd_sc_hd__a32o_1
X_9843_ clknet_leaf_35_i_clk rdata2\[27\] vssd1 vssd1 vccd1 vccd1 r_data2\[27\] sky130_fd_sc_hd__dfxtp_1
X_9774_ clknet_leaf_39_i_clk _0918_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6986_ _3349_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__clkbuf_1
X_5937_ reg_data\[24\]\[23\] _2453_ _2454_ reg_data\[28\]\[23\] _2516_ vssd1 vssd1
+ vccd1 vccd1 _2517_ sky130_fd_sc_hd__a221o_1
X_8725_ _4290_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__clkbuf_1
X_8656_ reg_data\[19\]\[1\] _3131_ _4252_ vssd1 vssd1 vccd1 vccd1 _4254_ sky130_fd_sc_hd__mux2_1
X_5868_ _1220_ vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__buf_2
X_7607_ _3210_ reg_data\[24\]\[4\] _3677_ vssd1 vssd1 vccd1 vccd1 _3682_ sky130_fd_sc_hd__mux2_1
X_5799_ reg_data\[6\]\[22\] _2207_ _2323_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__and3_1
X_8587_ _4217_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__clkbuf_1
X_4819_ reg_data\[4\]\[6\] _1074_ _1248_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__and3_1
X_7538_ reg_data\[23\]\[4\] _3137_ _3640_ vssd1 vssd1 vccd1 vccd1 _3645_ sky130_fd_sc_hd__mux2_1
X_7469_ _3210_ reg_data\[21\]\[4\] _3603_ vssd1 vssd1 vccd1 vccd1 _3608_ sky130_fd_sc_hd__mux2_1
X_9208_ clknet_leaf_9_i_clk _0352_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_9139_ clknet_leaf_17_i_clk _0283_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6840_ _3270_ vssd1 vssd1 vccd1 vccd1 _3271_ sky130_fd_sc_hd__buf_4
X_6771_ _3222_ reg_data\[22\]\[10\] _3223_ vssd1 vssd1 vccd1 vccd1 _3224_ sky130_fd_sc_hd__mux2_1
X_8510_ _3919_ reg_data\[18\]\[29\] _4166_ vssd1 vssd1 vccd1 vccd1 _4176_ sky130_fd_sc_hd__mux2_1
X_5722_ reg_data\[1\]\[20\] _1904_ _1905_ reg_data\[15\]\[20\] vssd1 vssd1 vccd1 vccd1
+ _2308_ sky130_fd_sc_hd__a22o_1
X_9490_ clknet_leaf_19_i_clk _0634_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_8441_ _4139_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__clkbuf_1
X_5653_ reg_data\[0\]\[19\] _1821_ _2238_ _2239_ _2240_ vssd1 vssd1 vccd1 vccd1 _2241_
+ sky130_fd_sc_hd__a2111o_1
X_8372_ _3917_ reg_data\[16\]\[28\] _4094_ vssd1 vssd1 vccd1 vccd1 _4103_ sky130_fd_sc_hd__mux2_1
X_5584_ reg_data\[25\]\[18\] _1810_ _2171_ _2172_ _2173_ vssd1 vssd1 vccd1 vccd1 _2174_
+ sky130_fd_sc_hd__a2111o_1
X_4604_ _1187_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__clkbuf_4
X_4535_ _0999_ _1155_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__and3_1
X_7323_ reg_data\[3\]\[0\] _3118_ _3529_ vssd1 vssd1 vccd1 vccd1 _3530_ sky130_fd_sc_hd__mux2_1
X_4466_ _1020_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__buf_4
X_7254_ _3492_ vssd1 vssd1 vccd1 vccd1 _3493_ sky130_fd_sc_hd__buf_4
X_6205_ reg_data\[2\]\[28\] _2443_ _2507_ _2508_ reg_data\[11\]\[28\] vssd1 vssd1
+ vccd1 vccd1 _2775_ sky130_fd_sc_hd__a32o_1
X_4397_ i_rs1[0] i_rs1[1] vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__nand2_1
X_7185_ _3455_ vssd1 vssd1 vccd1 vccd1 _3456_ sky130_fd_sc_hd__buf_4
X_6136_ reg_data\[25\]\[27\] _2416_ _2705_ _2706_ _2707_ vssd1 vssd1 vccd1 vccd1 _2708_
+ sky130_fd_sc_hd__a2111o_1
X_6067_ reg_data\[7\]\[26\] _2386_ _2639_ _2640_ _2641_ vssd1 vssd1 vccd1 vccd1 _2642_
+ sky130_fd_sc_hd__a2111o_1
X_5018_ reg_data\[25\]\[9\] _1141_ _1623_ _1624_ _1625_ vssd1 vssd1 vccd1 vccd1 _1626_
+ sky130_fd_sc_hd__a2111o_1
X_9826_ clknet_leaf_51_i_clk rdata2\[10\] vssd1 vssd1 vccd1 vccd1 r_data2\[10\] sky130_fd_sc_hd__dfxtp_1
X_6969_ _3260_ reg_data\[10\]\[28\] _3331_ vssd1 vssd1 vccd1 vccd1 _3340_ sky130_fd_sc_hd__mux2_1
X_9757_ clknet_leaf_0_i_clk _0901_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_8708_ reg_data\[19\]\[26\] _3183_ _4274_ vssd1 vssd1 vccd1 vccd1 _4281_ sky130_fd_sc_hd__mux2_1
X_9688_ clknet_leaf_61_i_clk _0832_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8639_ _4244_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_8990_ clknet_leaf_3_i_clk _0134_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_7941_ _3857_ reg_data\[9\]\[0\] _3859_ vssd1 vssd1 vccd1 vccd1 _3860_ sky130_fd_sc_hd__mux2_1
X_7872_ _3195_ reg_data\[28\]\[0\] _3822_ vssd1 vssd1 vccd1 vccd1 _3823_ sky130_fd_sc_hd__mux2_1
X_9611_ clknet_leaf_63_i_clk _0755_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6823_ _3258_ reg_data\[22\]\[27\] _3244_ vssd1 vssd1 vccd1 vccd1 _3259_ sky130_fd_sc_hd__mux2_1
X_6754_ i_data[5] vssd1 vssd1 vccd1 vccd1 _3212_ sky130_fd_sc_hd__clkbuf_4
X_9542_ clknet_leaf_45_i_clk _0686_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_5705_ reg_data\[18\]\[20\] _1816_ _2120_ vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__and3_1
X_9473_ clknet_leaf_5_i_clk _0617_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6685_ _3163_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__clkbuf_1
X_8424_ _3900_ reg_data\[17\]\[20\] _4130_ vssd1 vssd1 vccd1 vccd1 _4131_ sky130_fd_sc_hd__mux2_1
X_5636_ reg_data\[26\]\[19\] _1805_ _1806_ reg_data\[29\]\[19\] vssd1 vssd1 vccd1
+ vccd1 _2225_ sky130_fd_sc_hd__a22o_1
X_5567_ reg_data\[12\]\[18\] _1986_ _1606_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__and3_1
X_8355_ _4071_ vssd1 vssd1 vccd1 vccd1 _4094_ sky130_fd_sc_hd__buf_4
X_7306_ _3520_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__clkbuf_1
X_4518_ _1138_ _1139_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__and2_1
X_8286_ _4034_ vssd1 vssd1 vccd1 vccd1 _4057_ sky130_fd_sc_hd__buf_4
X_5498_ reg_data\[18\]\[17\] _1656_ _2090_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__and3_1
X_7237_ _3483_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__clkbuf_1
X_4449_ _1071_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__buf_2
X_7168_ reg_data\[7\]\[24\] _3179_ _3442_ vssd1 vssd1 vccd1 vccd1 _3447_ sky130_fd_sc_hd__mux2_1
X_7099_ _3252_ reg_data\[8\]\[24\] _3405_ vssd1 vssd1 vccd1 vccd1 _3410_ sky130_fd_sc_hd__mux2_1
X_6119_ reg_data\[12\]\[27\] _1082_ _2271_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__and3_1
X_9809_ clknet_leaf_35_i_clk rdata1\[25\] vssd1 vssd1 vccd1 vccd1 r_data1\[25\] sky130_fd_sc_hd__dfxtp_1
X_6470_ reg_data\[13\]\[1\] _1177_ _1190_ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__and3_1
X_5421_ reg_data\[12\]\[15\] _1960_ _2016_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__and3_1
X_5352_ reg_data\[3\]\[14\] _1815_ _1947_ _1948_ _1949_ vssd1 vssd1 vccd1 vccd1 _1950_
+ sky130_fd_sc_hd__a2111o_1
X_8140_ _3890_ reg_data\[13\]\[15\] _3974_ vssd1 vssd1 vccd1 vccd1 _3980_ sky130_fd_sc_hd__mux2_1
X_8071_ _3890_ reg_data\[30\]\[15\] _3937_ vssd1 vssd1 vccd1 vccd1 _3943_ sky130_fd_sc_hd__mux2_1
X_7022_ _3368_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__clkbuf_1
X_5283_ _1142_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__clkbuf_4
X_8973_ clknet_leaf_49_i_clk _0117_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_7924_ _3254_ reg_data\[28\]\[25\] _3844_ vssd1 vssd1 vccd1 vccd1 _3850_ sky130_fd_sc_hd__mux2_1
X_7855_ _3254_ reg_data\[27\]\[25\] _3807_ vssd1 vssd1 vccd1 vccd1 _3813_ sky130_fd_sc_hd__mux2_1
X_6806_ _3247_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__clkbuf_1
X_7786_ _3776_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__clkbuf_1
X_9525_ clknet_leaf_16_i_clk _0669_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_4998_ reg_data\[12\]\[9\] _1381_ _1606_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__and3_1
X_6737_ _3199_ vssd1 vssd1 vccd1 vccd1 _3200_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_63_i_clk clknet_3_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_9456_ clknet_leaf_31_i_clk _0600_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6668_ i_data[11] vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__buf_2
X_5619_ reg_data\[6\]\[19\] _2207_ _1716_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__and3_1
X_6599_ r_data2\[20\] _3105_ vssd1 vssd1 vccd1 vccd1 _3106_ sky130_fd_sc_hd__and2_1
X_9387_ clknet_leaf_57_i_clk _0531_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_8407_ _3884_ reg_data\[17\]\[12\] _4119_ vssd1 vssd1 vccd1 vccd1 _4122_ sky130_fd_sc_hd__mux2_1
X_8338_ _4085_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__clkbuf_1
X_8269_ _4048_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_16_i_clk clknet_3_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5970_ reg_data\[21\]\[24\] _2489_ _1943_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__and3_1
X_4921_ reg_data\[26\]\[7\] _1230_ _1232_ reg_data\[29\]\[7\] vssd1 vssd1 vccd1 vccd1
+ _1533_ sky130_fd_sc_hd__a22o_1
X_4852_ reg_data\[12\]\[6\] _1354_ _1226_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__and3_1
X_7640_ _3676_ vssd1 vssd1 vccd1 vccd1 _3699_ sky130_fd_sc_hd__buf_4
X_7571_ _3639_ vssd1 vssd1 vccd1 vccd1 _3662_ sky130_fd_sc_hd__clkbuf_4
X_4783_ reg_data\[25\]\[5\] _1141_ _1396_ _1397_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_
+ sky130_fd_sc_hd__a2111o_1
X_6522_ _3064_ vssd1 vssd1 vccd1 vccd1 o_data1[16] sky130_fd_sc_hd__buf_2
X_9310_ clknet_leaf_67_i_clk _0454_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_9241_ clknet_leaf_1_i_clk _0385_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6453_ reg_data\[8\]\[1\] _1115_ _1118_ reg_data\[10\]\[1\] _3013_ vssd1 vssd1 vccd1
+ vccd1 _3014_ sky130_fd_sc_hd__a221o_1
X_9172_ clknet_leaf_18_i_clk _0316_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_5404_ reg_data\[22\]\[15\] _1679_ _1622_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__and3_1
X_6384_ reg_data\[3\]\[0\] _1053_ _2944_ _2945_ _2946_ vssd1 vssd1 vccd1 vccd1 _2947_
+ sky130_fd_sc_hd__a2111o_1
X_8123_ _3873_ reg_data\[13\]\[7\] _3963_ vssd1 vssd1 vccd1 vccd1 _3971_ sky130_fd_sc_hd__mux2_1
X_5335_ reg_data\[2\]\[14\] _1613_ _1790_ _1791_ reg_data\[11\]\[14\] vssd1 vssd1
+ vccd1 vccd1 _1934_ sky130_fd_sc_hd__a32o_1
X_5266_ _1071_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__buf_2
X_8054_ _3873_ reg_data\[30\]\[7\] _3926_ vssd1 vssd1 vccd1 vccd1 _3934_ sky130_fd_sc_hd__mux2_1
X_7005_ _3359_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__clkbuf_1
X_5197_ _1122_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__buf_2
X_8956_ clknet_leaf_74_i_clk _0100_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_7907_ _3237_ reg_data\[28\]\[17\] _3833_ vssd1 vssd1 vccd1 vccd1 _3841_ sky130_fd_sc_hd__mux2_1
X_8887_ clknet_leaf_14_i_clk _0031_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_7838_ _3237_ reg_data\[27\]\[17\] _3796_ vssd1 vssd1 vccd1 vccd1 _3804_ sky130_fd_sc_hd__mux2_1
X_7769_ _3767_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__clkbuf_1
X_9508_ clknet_leaf_64_i_clk _0652_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_9439_ clknet_leaf_73_i_clk _0583_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5120_ reg_data\[7\]\[11\] _1081_ _1722_ _1723_ _1724_ vssd1 vssd1 vccd1 vccd1 _1725_
+ sky130_fd_sc_hd__a2111o_1
X_5051_ reg_data\[30\]\[10\] _1312_ _1313_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__and3_1
X_9790_ clknet_leaf_55_i_clk rdata1\[6\] vssd1 vssd1 vccd1 vccd1 r_data1\[6\] sky130_fd_sc_hd__dfxtp_1
X_8810_ _4323_ vssd1 vssd1 vccd1 vccd1 _4335_ sky130_fd_sc_hd__buf_4
X_8741_ _4298_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__clkbuf_1
X_5953_ reg_data\[0\]\[24\] _2381_ _2528_ _2529_ _2531_ vssd1 vssd1 vccd1 vccd1 _2532_
+ sky130_fd_sc_hd__a2111o_1
X_5884_ reg_data\[30\]\[23\] _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__and3_1
X_8672_ reg_data\[19\]\[9\] _3147_ _4252_ vssd1 vssd1 vccd1 vccd1 _4262_ sky130_fd_sc_hd__mux2_1
X_4904_ reg_data\[20\]\[7\] _1166_ _1180_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__and3_1
X_7623_ _3690_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__clkbuf_1
X_4835_ _1441_ _1445_ _1447_ _1449_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__or4_1
X_7554_ _3653_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__clkbuf_1
X_4766_ reg_data\[13\]\[5\] _1089_ _1257_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__and3_1
X_6505_ _3055_ vssd1 vssd1 vccd1 vccd1 o_data1[8] sky130_fd_sc_hd__buf_2
X_7485_ _3616_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__clkbuf_1
X_4697_ reg_data\[20\]\[4\] _1062_ _1315_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__and3_1
X_6436_ reg_data\[30\]\[1\] _2524_ _1056_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__and3_1
X_9224_ clknet_leaf_49_i_clk _0368_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6367_ reg_data\[23\]\[31\] _2440_ _2441_ reg_data\[19\]\[31\] vssd1 vssd1 vccd1
+ vccd1 _2931_ sky130_fd_sc_hd__a22o_1
X_9155_ clknet_leaf_63_i_clk _0299_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8106_ _3196_ _3124_ _3306_ vssd1 vssd1 vccd1 vccd1 _3961_ sky130_fd_sc_hd__and3_2
X_5318_ reg_data\[18\]\[14\] _1656_ _1483_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__and3_1
X_6298_ reg_data\[25\]\[30\] _2416_ _2861_ _2862_ _2863_ vssd1 vssd1 vccd1 vccd1 _2864_
+ sky130_fd_sc_hd__a2111o_1
X_9086_ clknet_leaf_2_i_clk _0230_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8037_ _3924_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__clkbuf_1
X_5249_ reg_data\[26\]\[12\] _1849_ _1850_ reg_data\[29\]\[12\] vssd1 vssd1 vccd1
+ vccd1 _1851_ sky130_fd_sc_hd__a22o_1
X_8939_ clknet_leaf_59_i_clk _0083_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_4620_ reg_data\[21\]\[3\] _1046_ _1240_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__and3_1
X_4551_ _1171_ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__and2_2
X_4482_ _1020_ _1094_ _1052_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__and3_4
X_7270_ _3501_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__clkbuf_1
X_6221_ reg_data\[3\]\[29\] _2376_ _2787_ _2788_ _2789_ vssd1 vssd1 vccd1 vccd1 _2790_
+ sky130_fd_sc_hd__a2111o_1
X_6152_ reg_data\[1\]\[27\] _2510_ _2511_ reg_data\[15\]\[27\] vssd1 vssd1 vccd1 vccd1
+ _2724_ sky130_fd_sc_hd__a22o_1
X_5103_ _1040_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__buf_4
X_6083_ reg_data\[18\]\[26\] _2422_ _2120_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__and3_1
X_9911_ clknet_leaf_40_i_clk _0981_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5034_ reg_data\[23\]\[9\] _1206_ _1209_ reg_data\[19\]\[9\] vssd1 vssd1 vccd1 vccd1
+ _1642_ sky130_fd_sc_hd__a22o_1
X_9842_ clknet_leaf_33_i_clk rdata2\[26\] vssd1 vssd1 vccd1 vccd1 r_data2\[26\] sky130_fd_sc_hd__dfxtp_1
X_9773_ clknet_leaf_40_i_clk _0917_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6985_ reg_data\[0\]\[3\] _3135_ _3345_ vssd1 vssd1 vccd1 vccd1 _3349_ sky130_fd_sc_hd__mux2_1
X_5936_ reg_data\[26\]\[23\] _2455_ _2456_ reg_data\[29\]\[23\] vssd1 vssd1 vccd1
+ vccd1 _2516_ sky130_fd_sc_hd__a22o_1
X_8724_ _3861_ reg_data\[29\]\[1\] _4288_ vssd1 vssd1 vccd1 vccd1 _4290_ sky130_fd_sc_hd__mux2_1
X_8655_ _4253_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__clkbuf_1
X_5867_ _1218_ vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__buf_2
X_7606_ _3681_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__clkbuf_1
X_5798_ _1069_ vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__clkbuf_4
X_8586_ _3857_ reg_data\[12\]\[0\] _4216_ vssd1 vssd1 vccd1 vccd1 _4217_ sky130_fd_sc_hd__mux2_1
X_4818_ reg_data\[6\]\[6\] _1072_ _1048_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__and3_1
X_4749_ _1366_ vssd1 vssd1 vccd1 vccd1 rdata2\[4\] sky130_fd_sc_hd__clkbuf_1
X_7537_ _3644_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__clkbuf_1
X_7468_ _3607_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__clkbuf_1
X_9207_ clknet_leaf_14_i_clk _0351_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6419_ reg_data\[7\]\[0\] _1184_ _2978_ _2979_ _2980_ vssd1 vssd1 vccd1 vccd1 _2981_
+ sky130_fd_sc_hd__a2111o_1
X_7399_ _3210_ reg_data\[20\]\[4\] _3565_ vssd1 vssd1 vccd1 vccd1 _3570_ sky130_fd_sc_hd__mux2_1
X_9138_ clknet_leaf_18_i_clk _0282_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_9069_ clknet_leaf_29_i_clk _0213_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6770_ _3201_ vssd1 vssd1 vccd1 vccd1 _3223_ sky130_fd_sc_hd__buf_4
X_5721_ reg_data\[2\]\[20\] _1837_ _1901_ _1902_ reg_data\[11\]\[20\] vssd1 vssd1
+ vccd1 vccd1 _2307_ sky130_fd_sc_hd__a32o_1
X_8440_ _3917_ reg_data\[17\]\[28\] _4130_ vssd1 vssd1 vccd1 vccd1 _4139_ sky130_fd_sc_hd__mux2_1
X_5652_ reg_data\[5\]\[19\] _1824_ _1954_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__and3_1
X_8371_ _4102_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__clkbuf_1
X_5583_ reg_data\[21\]\[18\] _2117_ _1510_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__and3_1
X_4603_ _1224_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__clkbuf_4
X_4534_ _0993_ _1006_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__nor2_2
X_7322_ _3528_ vssd1 vssd1 vccd1 vccd1 _3529_ sky130_fd_sc_hd__buf_4
X_7253_ _3125_ _3491_ vssd1 vssd1 vccd1 vccd1 _3492_ sky130_fd_sc_hd__nor2_2
X_4465_ reg_data\[13\]\[2\] _1085_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__and3_1
X_6204_ reg_data\[23\]\[28\] _2440_ _2441_ reg_data\[19\]\[28\] vssd1 vssd1 vccd1
+ vccd1 _2774_ sky130_fd_sc_hd__a22o_1
X_4396_ _1022_ vssd1 vssd1 vccd1 vccd1 rs1_mux\[4\] sky130_fd_sc_hd__clkinv_2
X_7184_ _3125_ _3268_ vssd1 vssd1 vccd1 vccd1 _3455_ sky130_fd_sc_hd__nor2_4
X_6135_ reg_data\[17\]\[27\] _1162_ _1148_ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__and3_1
X_6066_ reg_data\[13\]\[26\] _2214_ _2102_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__and3_1
X_5017_ reg_data\[17\]\[9\] _1509_ _1275_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__and3_1
X_9825_ clknet_leaf_54_i_clk rdata2\[9\] vssd1 vssd1 vccd1 vccd1 r_data2\[9\] sky130_fd_sc_hd__dfxtp_1
X_9756_ clknet_leaf_76_i_clk _0900_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6968_ _3339_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__clkbuf_1
X_8707_ _4280_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__clkbuf_1
X_5919_ reg_data\[5\]\[23\] _2430_ _1954_ vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__and3_1
X_6899_ reg_data\[2\]\[28\] _3187_ _3293_ vssd1 vssd1 vccd1 vccd1 _3302_ sky130_fd_sc_hd__mux2_1
X_9687_ clknet_leaf_14_i_clk _0831_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_8638_ _3911_ reg_data\[12\]\[25\] _4238_ vssd1 vssd1 vccd1 vccd1 _4244_ sky130_fd_sc_hd__mux2_1
X_8569_ _4207_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__clkbuf_1
X_7940_ _3858_ vssd1 vssd1 vccd1 vccd1 _3859_ sky130_fd_sc_hd__buf_4
X_7871_ _3821_ vssd1 vssd1 vccd1 vccd1 _3822_ sky130_fd_sc_hd__buf_4
X_6822_ i_data[27] vssd1 vssd1 vccd1 vccd1 _3258_ sky130_fd_sc_hd__clkbuf_4
X_9610_ clknet_leaf_51_i_clk _0754_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6753_ _3211_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__clkbuf_1
X_9541_ clknet_leaf_8_i_clk _0685_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5704_ reg_data\[25\]\[20\] _1810_ _2287_ _2288_ _2289_ vssd1 vssd1 vccd1 vccd1 _2290_
+ sky130_fd_sc_hd__a2111o_1
X_9472_ clknet_leaf_6_i_clk _0616_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6684_ reg_data\[4\]\[16\] _3162_ _3150_ vssd1 vssd1 vccd1 vccd1 _3163_ sky130_fd_sc_hd__mux2_1
X_8423_ _4107_ vssd1 vssd1 vccd1 vccd1 _4130_ sky130_fd_sc_hd__buf_4
X_5635_ reg_data\[8\]\[19\] _1797_ _1798_ reg_data\[10\]\[19\] _2223_ vssd1 vssd1
+ vccd1 vccd1 _2224_ sky130_fd_sc_hd__a221o_1
X_5566_ reg_data\[14\]\[18\] _1867_ _2156_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__and3_1
X_8354_ _4093_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__clkbuf_1
X_5497_ _1063_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__clkbuf_4
X_7305_ reg_data\[5\]\[24\] _3179_ _3515_ vssd1 vssd1 vccd1 vccd1 _3520_ sky130_fd_sc_hd__mux2_1
X_4517_ rs2_mux\[0\] _1006_ _1010_ rs2_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__and4_1
X_8285_ _4056_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__clkbuf_1
X_7236_ reg_data\[6\]\[24\] _3179_ _3478_ vssd1 vssd1 vccd1 vccd1 _3483_ sky130_fd_sc_hd__mux2_1
X_4448_ _1019_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__clkbuf_4
X_7167_ _3446_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__clkbuf_1
X_4379_ i_rs_valid rs2\[2\] vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__nor2_1
X_6118_ reg_data\[14\]\[27\] _2473_ _2156_ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__and3_1
X_7098_ _3409_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__clkbuf_1
X_6049_ reg_data\[24\]\[25\] _2453_ _2454_ reg_data\[28\]\[25\] _2624_ vssd1 vssd1
+ vccd1 vccd1 _2625_ sky130_fd_sc_hd__a221o_1
X_9808_ clknet_leaf_35_i_clk rdata1\[24\] vssd1 vssd1 vccd1 vccd1 r_data1\[24\] sky130_fd_sc_hd__dfxtp_1
X_9739_ clknet_leaf_26_i_clk _0883_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5420_ _1187_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__clkbuf_4
X_5351_ reg_data\[20\]\[14\] _1629_ _1743_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__and3_1
X_8070_ _3942_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__clkbuf_1
X_5282_ reg_data\[17\]\[13\] _1679_ _1147_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__and3_1
X_7021_ reg_data\[0\]\[20\] _3170_ _3367_ vssd1 vssd1 vccd1 vccd1 _3368_ sky130_fd_sc_hd__mux2_1
X_8972_ clknet_leaf_49_i_clk _0116_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_7923_ _3849_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__clkbuf_1
X_7854_ _3812_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__clkbuf_1
X_7785_ _3252_ reg_data\[26\]\[24\] _3771_ vssd1 vssd1 vccd1 vccd1 _3776_ sky130_fd_sc_hd__mux2_1
X_6805_ _3246_ reg_data\[22\]\[21\] _3244_ vssd1 vssd1 vccd1 vccd1 _3247_ sky130_fd_sc_hd__mux2_1
X_9524_ clknet_leaf_16_i_clk _0668_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_4997_ _1083_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__buf_2
X_6736_ i_rd[0] i_rd[1] i_write i_reset_n vssd1 vssd1 vccd1 vccd1 _3199_ sky130_fd_sc_hd__and4_1
X_9455_ clknet_leaf_32_i_clk _0599_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6667_ _3151_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__clkbuf_1
X_5618_ _1071_ vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__clkbuf_4
X_6598_ _3082_ vssd1 vssd1 vccd1 vccd1 _3105_ sky130_fd_sc_hd__clkbuf_2
X_9386_ clknet_leaf_55_i_clk _0530_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8406_ _4121_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__clkbuf_1
X_5549_ reg_data\[24\]\[17\] _1847_ _1848_ reg_data\[28\]\[17\] _2140_ vssd1 vssd1
+ vccd1 vccd1 _2141_ sky130_fd_sc_hd__a221o_1
X_8337_ _3882_ reg_data\[16\]\[11\] _4083_ vssd1 vssd1 vccd1 vccd1 _4085_ sky130_fd_sc_hd__mux2_1
X_8268_ _3882_ reg_data\[15\]\[11\] _4046_ vssd1 vssd1 vccd1 vccd1 _4048_ sky130_fd_sc_hd__mux2_1
X_8199_ _4011_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__clkbuf_1
X_7219_ reg_data\[6\]\[16\] _3162_ _3467_ vssd1 vssd1 vccd1 vccd1 _3474_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4920_ reg_data\[8\]\[7\] _1214_ _1217_ reg_data\[10\]\[7\] _1531_ vssd1 vssd1 vccd1
+ vccd1 _1532_ sky130_fd_sc_hd__a221o_1
X_4851_ reg_data\[14\]\[6\] _1189_ _1193_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__and3_1
X_7570_ _3661_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__clkbuf_1
X_4782_ reg_data\[22\]\[5\] _1150_ _1152_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__and3_1
X_6521_ r_data1\[16\] _3057_ vssd1 vssd1 vccd1 vccd1 _3064_ sky130_fd_sc_hd__and2_1
X_6452_ reg_data\[16\]\[1\] _1120_ _1122_ reg_data\[9\]\[1\] vssd1 vssd1 vccd1 vccd1
+ _3013_ sky130_fd_sc_hd__a22o_1
X_9240_ clknet_leaf_69_i_clk _0384_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_9171_ clknet_leaf_18_i_clk _0315_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5403_ _1999_ vssd1 vssd1 vccd1 vccd1 rdata1\[15\] sky130_fd_sc_hd__clkbuf_1
X_6383_ reg_data\[20\]\[0\] _1046_ _2035_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__and3_1
X_8122_ _3970_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__clkbuf_1
X_5334_ reg_data\[23\]\[14\] _1787_ _1788_ reg_data\[19\]\[14\] vssd1 vssd1 vccd1
+ vccd1 _1933_ sky130_fd_sc_hd__a22o_1
X_5265_ reg_data\[0\]\[13\] _1775_ _1862_ _1864_ _1865_ vssd1 vssd1 vccd1 vccd1 _1866_
+ sky130_fd_sc_hd__a2111o_1
X_8053_ _3933_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__clkbuf_1
X_5196_ _1120_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__clkbuf_4
X_7004_ reg_data\[0\]\[12\] _3154_ _3356_ vssd1 vssd1 vccd1 vccd1 _3359_ sky130_fd_sc_hd__mux2_1
X_8955_ clknet_leaf_71_i_clk _0099_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_8886_ clknet_leaf_16_i_clk _0030_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_7906_ _3840_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__clkbuf_1
X_7837_ _3803_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__clkbuf_1
X_7768_ _3235_ reg_data\[26\]\[16\] _3760_ vssd1 vssd1 vccd1 vccd1 _3767_ sky130_fd_sc_hd__mux2_1
X_6719_ _3186_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__clkbuf_1
X_7699_ _3730_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__clkbuf_1
X_9507_ clknet_leaf_7_i_clk _0651_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_9438_ clknet_leaf_73_i_clk _0582_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_9369_ clknet_leaf_67_i_clk _0513_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_5050_ reg_data\[18\]\[10\] _1656_ _1483_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_62_i_clk clknet_3_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5952_ reg_data\[5\]\[24\] _2097_ _2530_ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__and3_1
X_8740_ _3877_ reg_data\[29\]\[9\] _4288_ vssd1 vssd1 vccd1 vccd1 _4298_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_77_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4903_ reg_data\[30\]\[7\] _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__and3_1
X_5883_ reg_data\[18\]\[23\] _2261_ _2090_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__and3_1
X_8671_ _4261_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__clkbuf_1
X_7622_ _3225_ reg_data\[24\]\[11\] _3688_ vssd1 vssd1 vccd1 vccd1 _3690_ sky130_fd_sc_hd__mux2_1
X_4834_ reg_data\[24\]\[6\] _1127_ _1130_ reg_data\[28\]\[6\] _1448_ vssd1 vssd1 vccd1
+ vccd1 _1449_ sky130_fd_sc_hd__a221o_1
X_7553_ reg_data\[23\]\[11\] _3152_ _3651_ vssd1 vssd1 vccd1 vccd1 _3653_ sky130_fd_sc_hd__mux2_1
X_4765_ reg_data\[12\]\[5\] _1381_ _1128_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__and3_1
X_6504_ r_data1\[8\] _3046_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__and2_1
X_4696_ _1059_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__clkbuf_4
X_7484_ _3225_ reg_data\[21\]\[11\] _3614_ vssd1 vssd1 vccd1 vccd1 _3616_ sky130_fd_sc_hd__mux2_1
X_9223_ clknet_leaf_48_i_clk _0367_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[15\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_15_i_clk clknet_3_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_6435_ reg_data\[18\]\[1\] _1039_ _1063_ vssd1 vssd1 vccd1 vccd1 _2996_ sky130_fd_sc_hd__and3_1
X_6366_ _2917_ _2921_ _2925_ _2929_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__or4_4
X_9154_ clknet_leaf_68_i_clk _0298_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8105_ _3960_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__clkbuf_1
X_9085_ clknet_leaf_0_i_clk _0229_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_5317_ reg_data\[25\]\[14\] _1764_ _1913_ _1914_ _1915_ vssd1 vssd1 vccd1 vccd1 _1916_
+ sky130_fd_sc_hd__a2111o_1
X_6297_ reg_data\[17\]\[30\] _1162_ _1148_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__and3_1
X_8036_ _3923_ reg_data\[9\]\[31\] _3858_ vssd1 vssd1 vccd1 vccd1 _3924_ sky130_fd_sc_hd__mux2_1
X_5248_ _1231_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__clkbuf_4
X_5179_ reg_data\[12\]\[12\] _1381_ _1606_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__and3_1
X_8938_ clknet_leaf_56_i_clk _0082_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8869_ clknet_leaf_63_i_clk _0013_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_4550_ _0993_ _1006_ _1010_ _1013_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__and4_1
X_4481_ _1064_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__buf_4
X_6220_ reg_data\[30\]\[29\] _1046_ _1254_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__and3_1
X_6151_ reg_data\[2\]\[27\] _2443_ _2507_ _2508_ reg_data\[11\]\[27\] vssd1 vssd1
+ vccd1 vccd1 _2723_ sky130_fd_sc_hd__a32o_1
X_5102_ reg_data\[22\]\[11\] _1536_ _1651_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__and3_1
X_6082_ reg_data\[25\]\[26\] _2416_ _2653_ _2654_ _2655_ vssd1 vssd1 vccd1 vccd1 _2656_
+ sky130_fd_sc_hd__a2111o_1
X_5033_ _1626_ _1631_ _1636_ _1640_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__or4_1
X_9910_ clknet_leaf_49_i_clk _0980_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_9841_ clknet_leaf_35_i_clk rdata2\[25\] vssd1 vssd1 vccd1 vccd1 r_data2\[25\] sky130_fd_sc_hd__dfxtp_1
X_6984_ _3348_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__clkbuf_1
X_9772_ clknet_leaf_40_i_clk _0916_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5935_ reg_data\[8\]\[23\] _2447_ _2448_ reg_data\[10\]\[23\] _2514_ vssd1 vssd1
+ vccd1 vccd1 _2515_ sky130_fd_sc_hd__a221o_1
X_8723_ _4289_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__clkbuf_1
X_5866_ _1216_ vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__buf_2
X_8654_ reg_data\[19\]\[0\] _3118_ _4252_ vssd1 vssd1 vccd1 vccd1 _4253_ sky130_fd_sc_hd__mux2_1
X_7605_ _3208_ reg_data\[24\]\[3\] _3677_ vssd1 vssd1 vccd1 vccd1 _3681_ sky130_fd_sc_hd__mux2_1
X_4817_ reg_data\[3\]\[6\] _1054_ _1429_ _1430_ _1431_ vssd1 vssd1 vccd1 vccd1 _1432_
+ sky130_fd_sc_hd__a2111o_1
X_5797_ reg_data\[3\]\[22\] _2376_ _2377_ _2378_ _2379_ vssd1 vssd1 vccd1 vccd1 _2380_
+ sky130_fd_sc_hd__a2111o_1
X_8585_ _4215_ vssd1 vssd1 vccd1 vccd1 _4216_ sky130_fd_sc_hd__buf_4
X_4748_ _1357_ _1361_ _1363_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__or4_2
X_7536_ reg_data\[23\]\[3\] _3135_ _3640_ vssd1 vssd1 vccd1 vccd1 _3644_ sky130_fd_sc_hd__mux2_1
X_4679_ _1203_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__buf_4
X_7467_ _3208_ reg_data\[21\]\[3\] _3603_ vssd1 vssd1 vccd1 vccd1 _3607_ sky130_fd_sc_hd__mux2_1
X_9206_ clknet_leaf_20_i_clk _0350_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6418_ reg_data\[12\]\[0\] _2562_ _1289_ vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__and3_1
X_9137_ clknet_leaf_20_i_clk _0281_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_7398_ _3569_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__clkbuf_1
X_6349_ reg_data\[17\]\[31\] _1207_ _1147_ vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__and3_1
X_9068_ clknet_leaf_27_i_clk _0212_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8019_ _3912_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__clkbuf_1
X_5720_ reg_data\[23\]\[20\] _1834_ _1835_ reg_data\[19\]\[20\] vssd1 vssd1 vccd1
+ vccd1 _2306_ sky130_fd_sc_hd__a22o_1
X_5651_ reg_data\[4\]\[19\] _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__and3_1
X_8370_ _3915_ reg_data\[16\]\[27\] _4094_ vssd1 vssd1 vccd1 vccd1 _4102_ sky130_fd_sc_hd__mux2_1
X_4602_ _1166_ _1197_ _1212_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__and3_4
X_5582_ reg_data\[17\]\[18\] _1883_ _1395_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__and3_1
X_4533_ rs2_mux\[2\] rs2_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__nor2_1
X_7321_ _3269_ _3418_ vssd1 vssd1 vccd1 vccd1 _3528_ sky130_fd_sc_hd__nor2_4
X_7252_ _3126_ i_rd[0] i_rd[1] vssd1 vssd1 vccd1 vccd1 _3491_ sky130_fd_sc_hd__or3b_2
X_6203_ _2760_ _2764_ _2768_ _2772_ vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__or4_2
X_4464_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__clkbuf_4
X_4395_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__buf_6
X_7183_ _3454_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__clkbuf_1
X_6134_ reg_data\[21\]\[27\] _2489_ _1943_ vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__and3_1
X_6065_ reg_data\[12\]\[26\] _1082_ _2271_ vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__and3_1
X_5016_ reg_data\[21\]\[9\] _1272_ _1273_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__and3_1
X_9824_ clknet_leaf_55_i_clk rdata2\[8\] vssd1 vssd1 vccd1 vccd1 r_data2\[8\] sky130_fd_sc_hd__dfxtp_1
X_6967_ _3258_ reg_data\[10\]\[27\] _3331_ vssd1 vssd1 vccd1 vccd1 _3339_ sky130_fd_sc_hd__mux2_1
X_9755_ clknet_leaf_76_i_clk _0899_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_8706_ reg_data\[19\]\[25\] _3181_ _4274_ vssd1 vssd1 vccd1 vccd1 _4280_ sky130_fd_sc_hd__mux2_1
X_5918_ reg_data\[4\]\[23\] _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__and3_1
X_6898_ _3301_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__clkbuf_1
X_9686_ clknet_leaf_15_i_clk _0830_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_8637_ _4243_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__clkbuf_1
X_5849_ reg_data\[5\]\[22\] _2430_ _1954_ vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__and3_1
X_8568_ reg_data\[1\]\[24\] _3179_ _4202_ vssd1 vssd1 vccd1 vccd1 _4207_ sky130_fd_sc_hd__mux2_1
X_7519_ _3260_ reg_data\[21\]\[28\] _3625_ vssd1 vssd1 vccd1 vccd1 _3634_ sky130_fd_sc_hd__mux2_1
X_8499_ _4170_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__clkbuf_1
X_7870_ _3127_ _3820_ vssd1 vssd1 vccd1 vccd1 _3821_ sky130_fd_sc_hd__or2_4
X_6821_ _3257_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__clkbuf_1
X_9540_ clknet_leaf_65_i_clk _0684_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_6752_ _3210_ reg_data\[22\]\[4\] _3202_ vssd1 vssd1 vccd1 vccd1 _3211_ sky130_fd_sc_hd__mux2_1
X_5703_ reg_data\[21\]\[20\] _2117_ _1510_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__and3_1
X_6683_ i_data[16] vssd1 vssd1 vccd1 vccd1 _3162_ sky130_fd_sc_hd__clkbuf_4
X_9471_ clknet_leaf_3_i_clk _0615_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8422_ _4129_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__clkbuf_1
X_5634_ reg_data\[16\]\[19\] _1799_ _1800_ reg_data\[9\]\[19\] vssd1 vssd1 vccd1 vccd1
+ _2223_ sky130_fd_sc_hd__a22o_1
X_8353_ _3898_ reg_data\[16\]\[19\] _4083_ vssd1 vssd1 vccd1 vccd1 _4093_ sky130_fd_sc_hd__mux2_1
X_7304_ _3519_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__clkbuf_1
X_5565_ _1056_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__clkbuf_4
X_4516_ _0997_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__buf_2
X_5496_ reg_data\[25\]\[17\] _1764_ _2084_ _2085_ _2088_ vssd1 vssd1 vccd1 vccd1 _2089_
+ sky130_fd_sc_hd__a2111o_1
X_8284_ _3898_ reg_data\[15\]\[19\] _4046_ vssd1 vssd1 vccd1 vccd1 _4056_ sky130_fd_sc_hd__mux2_1
X_7235_ _3482_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__clkbuf_1
X_4447_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__clkbuf_4
X_7166_ reg_data\[7\]\[23\] _3177_ _3442_ vssd1 vssd1 vccd1 vccd1 _3446_ sky130_fd_sc_hd__mux2_1
X_6117_ reg_data\[0\]\[27\] _2381_ _2687_ _2688_ _2689_ vssd1 vssd1 vccd1 vccd1 _2690_
+ sky130_fd_sc_hd__a2111o_1
X_4378_ i_rs2[0] i_rs2[1] i_rs2[2] vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__o21ai_1
X_7097_ _3250_ reg_data\[8\]\[23\] _3405_ vssd1 vssd1 vccd1 vccd1 _3409_ sky130_fd_sc_hd__mux2_1
X_6048_ reg_data\[26\]\[25\] _2455_ _2456_ reg_data\[29\]\[25\] vssd1 vssd1 vccd1
+ vccd1 _2624_ sky130_fd_sc_hd__a22o_1
X_9807_ clknet_leaf_36_i_clk rdata1\[23\] vssd1 vssd1 vccd1 vccd1 r_data1\[23\] sky130_fd_sc_hd__dfxtp_1
X_7999_ _3898_ reg_data\[9\]\[19\] _3880_ vssd1 vssd1 vccd1 vccd1 _3899_ sky130_fd_sc_hd__mux2_1
X_9738_ clknet_leaf_26_i_clk _0882_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_9669_ clknet_leaf_45_i_clk _0813_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5350_ reg_data\[30\]\[14\] _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__and3_1
X_5281_ _1881_ vssd1 vssd1 vccd1 vccd1 rdata1\[13\] sky130_fd_sc_hd__clkbuf_1
X_7020_ _3344_ vssd1 vssd1 vccd1 vccd1 _3367_ sky130_fd_sc_hd__buf_4
X_8971_ clknet_leaf_52_i_clk _0115_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_7922_ _3252_ reg_data\[28\]\[24\] _3844_ vssd1 vssd1 vccd1 vccd1 _3849_ sky130_fd_sc_hd__mux2_1
X_7853_ _3252_ reg_data\[27\]\[24\] _3807_ vssd1 vssd1 vccd1 vccd1 _3812_ sky130_fd_sc_hd__mux2_1
X_7784_ _3775_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__clkbuf_1
X_6804_ i_data[21] vssd1 vssd1 vccd1 vccd1 _3246_ sky130_fd_sc_hd__buf_2
X_4996_ reg_data\[14\]\[9\] _1253_ _1379_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__and3_1
X_9523_ clknet_leaf_18_i_clk _0667_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6735_ i_rd[4] _3196_ _3197_ vssd1 vssd1 vccd1 vccd1 _3198_ sky130_fd_sc_hd__and3_2
X_9454_ clknet_leaf_32_i_clk _0598_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6666_ reg_data\[4\]\[10\] _3149_ _3150_ vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__mux2_1
X_6597_ _3104_ vssd1 vssd1 vccd1 vccd1 o_data2[19] sky130_fd_sc_hd__buf_2
X_5617_ reg_data\[3\]\[19\] _1770_ _2202_ _2203_ _2205_ vssd1 vssd1 vccd1 vccd1 _2206_
+ sky130_fd_sc_hd__a2111o_1
X_9385_ clknet_leaf_57_i_clk _0529_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_8405_ _3882_ reg_data\[17\]\[11\] _4119_ vssd1 vssd1 vccd1 vccd1 _4121_ sky130_fd_sc_hd__mux2_1
X_5548_ reg_data\[26\]\[17\] _1849_ _1850_ reg_data\[29\]\[17\] vssd1 vssd1 vccd1
+ vccd1 _2140_ sky130_fd_sc_hd__a22o_1
X_8336_ _4084_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__clkbuf_1
X_8267_ _4047_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__clkbuf_1
X_7218_ _3473_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
X_5479_ reg_data\[7\]\[16\] _1827_ _2070_ _2071_ _2072_ vssd1 vssd1 vccd1 vccd1 _2073_
+ sky130_fd_sc_hd__a2111o_1
X_8198_ _3879_ reg_data\[14\]\[10\] _4010_ vssd1 vssd1 vccd1 vccd1 _4011_ sky130_fd_sc_hd__mux2_1
X_7149_ reg_data\[7\]\[15\] _3160_ _3431_ vssd1 vssd1 vccd1 vccd1 _3437_ sky130_fd_sc_hd__mux2_1
X_4850_ reg_data\[13\]\[6\] _1186_ _1191_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__and3_1
X_6520_ _3063_ vssd1 vssd1 vccd1 vccd1 o_data1[15] sky130_fd_sc_hd__buf_2
X_4781_ reg_data\[21\]\[5\] _1272_ _1273_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__and3_1
X_6451_ reg_data\[27\]\[1\] _1095_ _3009_ _3010_ _3011_ vssd1 vssd1 vccd1 vccd1 _3012_
+ sky130_fd_sc_hd__a2111o_1
X_9170_ clknet_leaf_19_i_clk _0314_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6382_ reg_data\[30\]\[0\] _2524_ _1056_ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__and3_1
X_5402_ _1990_ _1994_ _1996_ _1998_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__or4_1
X_5333_ _1916_ _1922_ _1927_ _1931_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__or4_1
X_8121_ _3871_ reg_data\[13\]\[6\] _3963_ vssd1 vssd1 vccd1 vccd1 _3970_ sky130_fd_sc_hd__mux2_1
X_5264_ reg_data\[5\]\[13\] _1490_ _1250_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__and3_1
X_8052_ _3871_ reg_data\[30\]\[6\] _3926_ vssd1 vssd1 vccd1 vccd1 _3933_ sky130_fd_sc_hd__mux2_1
X_7003_ _3358_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__clkbuf_1
X_5195_ _1118_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__clkbuf_4
X_8954_ clknet_leaf_61_i_clk _0098_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8885_ clknet_leaf_16_i_clk _0029_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_7905_ _3235_ reg_data\[28\]\[16\] _3833_ vssd1 vssd1 vccd1 vccd1 _3840_ sky130_fd_sc_hd__mux2_1
X_7836_ _3235_ reg_data\[27\]\[16\] _3796_ vssd1 vssd1 vccd1 vccd1 _3803_ sky130_fd_sc_hd__mux2_1
X_4979_ reg_data\[24\]\[8\] _1225_ _1228_ reg_data\[28\]\[8\] _1588_ vssd1 vssd1 vccd1
+ vccd1 _1589_ sky130_fd_sc_hd__a221o_1
X_7767_ _3766_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__clkbuf_1
X_6718_ reg_data\[4\]\[27\] _3185_ _3171_ vssd1 vssd1 vccd1 vccd1 _3186_ sky130_fd_sc_hd__mux2_1
X_7698_ _3233_ reg_data\[25\]\[15\] _3724_ vssd1 vssd1 vccd1 vccd1 _3730_ sky130_fd_sc_hd__mux2_1
X_9506_ clknet_leaf_7_i_clk _0650_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_9437_ clknet_leaf_71_i_clk _0581_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6649_ i_data[5] vssd1 vssd1 vccd1 vccd1 _3139_ sky130_fd_sc_hd__buf_2
X_9368_ clknet_leaf_61_i_clk _0512_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_9299_ clknet_leaf_35_i_clk _0443_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_8319_ _4075_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__clkbuf_1
X_5951_ _1043_ vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__buf_2
X_8670_ reg_data\[19\]\[8\] _3145_ _4252_ vssd1 vssd1 vccd1 vccd1 _4261_ sky130_fd_sc_hd__mux2_1
X_4902_ reg_data\[18\]\[7\] _1159_ _1513_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__and3_1
X_5882_ reg_data\[25\]\[23\] _2370_ _2460_ _2461_ _2462_ vssd1 vssd1 vccd1 vccd1 _2463_
+ sky130_fd_sc_hd__a2111o_1
X_4833_ reg_data\[26\]\[6\] _1132_ _1134_ reg_data\[29\]\[6\] vssd1 vssd1 vccd1 vccd1
+ _1448_ sky130_fd_sc_hd__a22o_1
X_7621_ _3689_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__clkbuf_1
X_7552_ _3652_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__clkbuf_1
X_4764_ _1067_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__buf_2
X_6503_ _3054_ vssd1 vssd1 vccd1 vccd1 o_data1[7] sky130_fd_sc_hd__buf_2
X_7483_ _3615_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__clkbuf_1
X_6434_ reg_data\[25\]\[1\] _1036_ _2992_ _2993_ _2994_ vssd1 vssd1 vccd1 vccd1 _2995_
+ sky130_fd_sc_hd__a2111o_1
X_9222_ clknet_leaf_49_i_clk _0366_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_4695_ reg_data\[30\]\[4\] _1312_ _1313_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__and3_1
X_6365_ reg_data\[7\]\[31\] _2433_ _2926_ _2927_ _2928_ vssd1 vssd1 vccd1 vccd1 _2929_
+ sky130_fd_sc_hd__a2111o_1
X_9153_ clknet_leaf_5_i_clk _0297_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6296_ reg_data\[21\]\[30\] _2489_ _1943_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__and3_1
X_8104_ _3923_ reg_data\[30\]\[31\] _3925_ vssd1 vssd1 vccd1 vccd1 _3960_ sky130_fd_sc_hd__mux2_1
X_5316_ reg_data\[17\]\[14\] _1480_ _1108_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__and3_1
X_9084_ clknet_leaf_5_i_clk _0228_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_8035_ i_data[31] vssd1 vssd1 vccd1 vccd1 _3923_ sky130_fd_sc_hd__clkbuf_4
X_5247_ _1229_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__clkbuf_4
X_5178_ reg_data\[14\]\[12\] _1253_ _1379_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__and3_1
X_8937_ clknet_leaf_56_i_clk _0081_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_8868_ clknet_leaf_63_i_clk _0012_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_7819_ _3218_ reg_data\[27\]\[8\] _3785_ vssd1 vssd1 vccd1 vccd1 _3794_ sky130_fd_sc_hd__mux2_1
X_8799_ _4329_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__clkbuf_1
X_4480_ _1021_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__buf_4
X_6150_ reg_data\[23\]\[27\] _2440_ _2441_ reg_data\[19\]\[27\] vssd1 vssd1 vccd1
+ vccd1 _2722_ sky130_fd_sc_hd__a22o_1
X_5101_ _1706_ vssd1 vssd1 vccd1 vccd1 rdata2\[10\] sky130_fd_sc_hd__dlymetal6s2s_1
X_6081_ reg_data\[21\]\[26\] _2117_ _1510_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__and3_1
X_5032_ reg_data\[7\]\[9\] _1185_ _1637_ _1638_ _1639_ vssd1 vssd1 vccd1 vccd1 _1640_
+ sky130_fd_sc_hd__a2111o_1
X_9840_ clknet_leaf_33_i_clk rdata2\[24\] vssd1 vssd1 vccd1 vccd1 r_data2\[24\] sky130_fd_sc_hd__dfxtp_1
X_6983_ reg_data\[0\]\[2\] _3133_ _3345_ vssd1 vssd1 vccd1 vccd1 _3348_ sky130_fd_sc_hd__mux2_1
X_9771_ clknet_leaf_59_i_clk _0915_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5934_ reg_data\[16\]\[23\] _2449_ _2450_ reg_data\[9\]\[23\] vssd1 vssd1 vccd1 vccd1
+ _2514_ sky130_fd_sc_hd__a22o_1
X_8722_ _3857_ reg_data\[29\]\[0\] _4288_ vssd1 vssd1 vccd1 vccd1 _4289_ sky130_fd_sc_hd__mux2_1
X_5865_ _1213_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__buf_2
X_8653_ _4251_ vssd1 vssd1 vccd1 vccd1 _4252_ sky130_fd_sc_hd__buf_4
X_7604_ _3680_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__clkbuf_1
X_4816_ reg_data\[30\]\[6\] _1062_ _1254_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__and3_1
X_5796_ reg_data\[30\]\[22\] _2204_ _1254_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__and3_1
X_8584_ _3381_ _3961_ vssd1 vssd1 vccd1 vccd1 _4215_ sky130_fd_sc_hd__nand2_2
X_4747_ reg_data\[24\]\[4\] _1225_ _1228_ reg_data\[28\]\[4\] _1364_ vssd1 vssd1 vccd1
+ vccd1 _1365_ sky130_fd_sc_hd__a221o_1
X_7535_ _3643_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__clkbuf_1
X_4678_ _1202_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__buf_4
X_7466_ _3606_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__clkbuf_1
X_9205_ clknet_leaf_20_i_clk _0349_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6417_ reg_data\[14\]\[0\] _1186_ _1344_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__and3_1
X_7397_ _3208_ reg_data\[20\]\[3\] _3565_ vssd1 vssd1 vccd1 vccd1 _3569_ sky130_fd_sc_hd__mux2_1
X_9136_ clknet_leaf_20_i_clk _0280_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6348_ _2912_ vssd1 vssd1 vccd1 vccd1 rdata1\[31\] sky130_fd_sc_hd__clkbuf_1
X_6279_ reg_data\[0\]\[30\] _2381_ _2843_ _2844_ _2845_ vssd1 vssd1 vccd1 vccd1 _2846_
+ sky130_fd_sc_hd__a2111o_1
X_9067_ clknet_leaf_27_i_clk _0211_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_8018_ _3911_ reg_data\[9\]\[25\] _3901_ vssd1 vssd1 vccd1 vccd1 _3912_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_61_i_clk clknet_3_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_76_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_14_i_clk clknet_3_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5650_ reg_data\[6\]\[19\] _1951_ _2237_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__and3_1
X_4601_ reg_data\[8\]\[2\] _1214_ _1217_ reg_data\[10\]\[2\] _1222_ vssd1 vssd1 vccd1
+ vccd1 _1223_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_29_i_clk clknet_3_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5581_ reg_data\[22\]\[18\] _1679_ _1622_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__and3_1
X_7320_ _3527_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__clkbuf_1
X_4532_ reg_data\[25\]\[2\] _1141_ _1145_ _1149_ _1153_ vssd1 vssd1 vccd1 vccd1 _1154_
+ sky130_fd_sc_hd__a2111o_1
X_4463_ rs1_mux\[0\] _1026_ rs1_mux\[2\] rs1_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1086_
+ sky130_fd_sc_hd__and4_2
X_7251_ _3490_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__clkbuf_1
X_6202_ reg_data\[7\]\[28\] _2433_ _2769_ _2770_ _2771_ vssd1 vssd1 vccd1 vccd1 _2772_
+ sky130_fd_sc_hd__a2111o_1
X_7182_ reg_data\[7\]\[31\] _3193_ _3419_ vssd1 vssd1 vccd1 vccd1 _3454_ sky130_fd_sc_hd__mux2_1
X_4394_ _1020_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__buf_6
X_6133_ reg_data\[22\]\[27\] _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__and3_1
X_6064_ reg_data\[14\]\[26\] _2473_ _2156_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__and3_1
X_5015_ reg_data\[22\]\[9\] _1143_ _1622_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__and3_1
X_9823_ clknet_leaf_72_i_clk rdata2\[7\] vssd1 vssd1 vccd1 vccd1 r_data2\[7\] sky130_fd_sc_hd__dfxtp_2
X_6966_ _3338_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__clkbuf_1
X_9754_ clknet_leaf_74_i_clk _0898_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8705_ _4279_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__clkbuf_1
X_5917_ reg_data\[6\]\[23\] _1951_ _2237_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__and3_1
X_6897_ reg_data\[2\]\[27\] _3185_ _3293_ vssd1 vssd1 vccd1 vccd1 _3301_ sky130_fd_sc_hd__mux2_1
X_9685_ clknet_leaf_16_i_clk _0829_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_8636_ _3909_ reg_data\[12\]\[24\] _4238_ vssd1 vssd1 vccd1 vccd1 _4243_ sky130_fd_sc_hd__mux2_1
X_5848_ _1171_ vssd1 vssd1 vccd1 vccd1 _2430_ sky130_fd_sc_hd__buf_2
X_8567_ _4206_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__clkbuf_1
X_5779_ reg_data\[1\]\[21\] _1904_ _1905_ reg_data\[15\]\[21\] vssd1 vssd1 vccd1 vccd1
+ _2363_ sky130_fd_sc_hd__a22o_1
X_7518_ _3633_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__clkbuf_1
X_8498_ _3907_ reg_data\[18\]\[23\] _4166_ vssd1 vssd1 vccd1 vccd1 _4170_ sky130_fd_sc_hd__mux2_1
X_7449_ _3260_ reg_data\[20\]\[28\] _3587_ vssd1 vssd1 vccd1 vccd1 _3596_ sky130_fd_sc_hd__mux2_1
X_9119_ clknet_leaf_3_i_clk _0263_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6820_ _3256_ reg_data\[22\]\[26\] _3244_ vssd1 vssd1 vccd1 vccd1 _3257_ sky130_fd_sc_hd__mux2_1
X_6751_ i_data[4] vssd1 vssd1 vccd1 vccd1 _3210_ sky130_fd_sc_hd__clkbuf_4
X_5702_ reg_data\[17\]\[20\] _1883_ _1395_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__and3_1
X_9470_ clknet_leaf_3_i_clk _0614_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6682_ _3161_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__clkbuf_1
X_8421_ _3898_ reg_data\[17\]\[19\] _4119_ vssd1 vssd1 vccd1 vccd1 _4129_ sky130_fd_sc_hd__mux2_1
X_5633_ reg_data\[27\]\[19\] _1786_ _2218_ _2220_ _2221_ vssd1 vssd1 vccd1 vccd1 _2222_
+ sky130_fd_sc_hd__a2111o_1
X_5564_ reg_data\[0\]\[18\] _1775_ _2152_ _2153_ _2154_ vssd1 vssd1 vccd1 vccd1 _2155_
+ sky130_fd_sc_hd__a2111o_1
X_8352_ _4092_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__clkbuf_1
X_7303_ reg_data\[5\]\[23\] _3177_ _3515_ vssd1 vssd1 vccd1 vccd1 _3519_ sky130_fd_sc_hd__mux2_1
X_4515_ _1137_ vssd1 vssd1 vccd1 vccd1 rdata1\[2\] sky130_fd_sc_hd__dlymetal6s2s_1
X_5495_ reg_data\[21\]\[17\] _2086_ _2087_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__and3_1
X_8283_ _4055_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__clkbuf_1
X_7234_ reg_data\[6\]\[23\] _3177_ _3478_ vssd1 vssd1 vccd1 vccd1 _3482_ sky130_fd_sc_hd__mux2_1
X_4446_ _1067_ _1068_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__and2_1
X_7165_ _3445_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__clkbuf_1
X_4377_ i_rs2[0] i_rs2[2] i_rs2[1] vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__or3_1
X_6116_ reg_data\[5\]\[27\] _1085_ _2530_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__and3_1
X_7096_ _3408_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__clkbuf_1
X_6047_ reg_data\[8\]\[25\] _2447_ _2448_ reg_data\[10\]\[25\] _2622_ vssd1 vssd1
+ vccd1 vccd1 _2623_ sky130_fd_sc_hd__a221o_1
X_9806_ clknet_leaf_39_i_clk rdata1\[22\] vssd1 vssd1 vccd1 vccd1 r_data1\[22\] sky130_fd_sc_hd__dfxtp_1
X_7998_ i_data[19] vssd1 vssd1 vccd1 vccd1 _3898_ sky130_fd_sc_hd__clkbuf_4
X_9737_ clknet_leaf_26_i_clk _0881_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6949_ _3329_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__clkbuf_1
X_9668_ clknet_leaf_47_i_clk _0812_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8619_ _3892_ reg_data\[12\]\[16\] _4227_ vssd1 vssd1 vccd1 vccd1 _4234_ sky130_fd_sc_hd__mux2_1
X_9599_ clknet_leaf_72_i_clk _0743_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5280_ _1872_ _1876_ _1878_ _1880_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__or4_1
X_8970_ clknet_leaf_50_i_clk _0114_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_7921_ _3848_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__clkbuf_1
X_7852_ _3811_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__clkbuf_1
X_7783_ _3250_ reg_data\[26\]\[23\] _3771_ vssd1 vssd1 vccd1 vccd1 _3775_ sky130_fd_sc_hd__mux2_1
X_6803_ _3245_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__clkbuf_1
X_4995_ reg_data\[0\]\[9\] _1070_ _1601_ _1602_ _1603_ vssd1 vssd1 vccd1 vccd1 _1604_
+ sky130_fd_sc_hd__a2111o_1
X_9522_ clknet_leaf_17_i_clk _0666_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6734_ _3122_ _3123_ vssd1 vssd1 vccd1 vccd1 _3197_ sky130_fd_sc_hd__and2_1
X_9453_ clknet_leaf_50_i_clk _0597_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6665_ _3128_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__buf_6
X_8404_ _4120_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__clkbuf_1
X_5616_ reg_data\[30\]\[19\] _2204_ _1254_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__and3_1
X_9384_ clknet_leaf_55_i_clk _0528_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6596_ r_data2\[19\] _3094_ vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__and2_1
X_8335_ _3879_ reg_data\[16\]\[10\] _4083_ vssd1 vssd1 vccd1 vccd1 _4084_ sky130_fd_sc_hd__mux2_1
X_5547_ reg_data\[8\]\[17\] _1841_ _1842_ reg_data\[10\]\[17\] _2138_ vssd1 vssd1
+ vccd1 vccd1 _2139_ sky130_fd_sc_hd__a221o_1
X_8266_ _3879_ reg_data\[15\]\[10\] _4046_ vssd1 vssd1 vccd1 vccd1 _4047_ sky130_fd_sc_hd__mux2_1
X_5478_ reg_data\[12\]\[16\] _1960_ _2016_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__and3_1
X_4429_ _1015_ _1026_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__nor2_2
X_7217_ reg_data\[6\]\[15\] _3160_ _3467_ vssd1 vssd1 vccd1 vccd1 _3473_ sky130_fd_sc_hd__mux2_1
X_8197_ _3998_ vssd1 vssd1 vccd1 vccd1 _4010_ sky130_fd_sc_hd__buf_4
X_7148_ _3436_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__clkbuf_1
X_7079_ _3399_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_1
X_4780_ reg_data\[17\]\[5\] _1143_ _1395_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__and3_1
X_6450_ reg_data\[1\]\[1\] _1103_ _1108_ _1110_ reg_data\[15\]\[1\] vssd1 vssd1 vccd1
+ vccd1 _3011_ sky130_fd_sc_hd__a32o_1
X_6381_ reg_data\[18\]\[0\] _1039_ _1063_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__and3_1
X_5401_ reg_data\[24\]\[15\] _1803_ _1804_ reg_data\[28\]\[15\] _1997_ vssd1 vssd1
+ vccd1 vccd1 _1998_ sky130_fd_sc_hd__a221o_1
X_8120_ _3969_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__clkbuf_1
X_5332_ reg_data\[7\]\[14\] _1780_ _1928_ _1929_ _1930_ vssd1 vssd1 vccd1 vccd1 _1931_
+ sky130_fd_sc_hd__a2111o_1
X_5263_ reg_data\[4\]\[13\] _1718_ _1863_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__and3_1
X_8051_ _3932_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__clkbuf_1
X_7002_ reg_data\[0\]\[11\] _3152_ _3356_ vssd1 vssd1 vccd1 vccd1 _3358_ sky130_fd_sc_hd__mux2_1
X_5194_ _1115_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__clkbuf_4
X_8953_ clknet_leaf_67_i_clk _0097_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8884_ clknet_leaf_16_i_clk _0028_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_7904_ _3839_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__clkbuf_1
X_7835_ _3802_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__clkbuf_1
X_4978_ reg_data\[26\]\[8\] _1230_ _1232_ reg_data\[29\]\[8\] vssd1 vssd1 vccd1 vccd1
+ _1588_ sky130_fd_sc_hd__a22o_1
X_7766_ _3233_ reg_data\[26\]\[15\] _3760_ vssd1 vssd1 vccd1 vccd1 _3766_ sky130_fd_sc_hd__mux2_1
X_9505_ clknet_leaf_7_i_clk _0649_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6717_ i_data[27] vssd1 vssd1 vccd1 vccd1 _3185_ sky130_fd_sc_hd__buf_4
X_7697_ _3729_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__clkbuf_1
X_9436_ clknet_leaf_74_i_clk _0580_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6648_ _3138_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__clkbuf_1
X_9367_ clknet_leaf_38_i_clk _0511_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_8318_ _3863_ reg_data\[16\]\[2\] _4072_ vssd1 vssd1 vccd1 vccd1 _4075_ sky130_fd_sc_hd__mux2_1
X_6579_ _3095_ vssd1 vssd1 vccd1 vccd1 o_data2[10] sky130_fd_sc_hd__buf_2
X_9298_ clknet_leaf_34_i_clk _0442_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_8249_ _3863_ reg_data\[15\]\[2\] _4035_ vssd1 vssd1 vccd1 vccd1 _4038_ sky130_fd_sc_hd__mux2_1
X_5950_ reg_data\[4\]\[24\] _2325_ _2469_ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__and3_1
X_4901_ _1167_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__clkbuf_4
X_5881_ reg_data\[17\]\[23\] _2086_ _1238_ vssd1 vssd1 vccd1 vccd1 _2462_ sky130_fd_sc_hd__and3_1
X_7620_ _3222_ reg_data\[24\]\[10\] _3688_ vssd1 vssd1 vccd1 vccd1 _3689_ sky130_fd_sc_hd__mux2_1
X_4832_ reg_data\[8\]\[6\] _1116_ _1119_ reg_data\[10\]\[6\] _1446_ vssd1 vssd1 vccd1
+ vccd1 _1447_ sky130_fd_sc_hd__a221o_1
X_7551_ reg_data\[23\]\[10\] _3149_ _3651_ vssd1 vssd1 vccd1 vccd1 _3652_ sky130_fd_sc_hd__mux2_1
X_4763_ reg_data\[14\]\[5\] _1253_ _1379_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__and3_1
X_4694_ _1056_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__clkbuf_4
X_6502_ r_data1\[7\] _3046_ vssd1 vssd1 vccd1 vccd1 _3054_ sky130_fd_sc_hd__and2_1
X_7482_ _3222_ reg_data\[21\]\[10\] _3614_ vssd1 vssd1 vccd1 vccd1 _3615_ sky130_fd_sc_hd__mux2_1
X_6433_ reg_data\[21\]\[1\] _1058_ _1044_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__and3_1
X_9221_ clknet_leaf_64_i_clk _0365_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6364_ reg_data\[12\]\[31\] _2562_ _1289_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__and3_1
X_9152_ clknet_leaf_3_i_clk _0296_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6295_ reg_data\[22\]\[30\] _1207_ _1151_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__and3_1
X_8103_ _3959_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__clkbuf_1
X_9083_ clknet_leaf_3_i_clk _0227_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5315_ reg_data\[21\]\[14\] _1766_ _1044_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__and3_1
X_8034_ _3922_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__clkbuf_1
X_5246_ _1227_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__clkbuf_4
X_5177_ _1080_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__clkbuf_4
X_8936_ clknet_leaf_56_i_clk _0080_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_8867_ clknet_leaf_63_i_clk _0011_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8798_ reg_data\[11\]\[4\] i_data[4] _4324_ vssd1 vssd1 vccd1 vccd1 _4329_ sky130_fd_sc_hd__mux2_1
X_7818_ _3793_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__clkbuf_1
X_7749_ _3216_ reg_data\[26\]\[7\] _3749_ vssd1 vssd1 vccd1 vccd1 _3757_ sky130_fd_sc_hd__mux2_1
X_9419_ clknet_leaf_59_i_clk _0563_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6080_ reg_data\[17\]\[26\] _2489_ _1395_ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__and3_1
X_5100_ _1697_ _1701_ _1703_ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__or4_1
X_5031_ reg_data\[12\]\[9\] _1354_ _1226_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__and3_1
X_9770_ clknet_leaf_56_i_clk _0914_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6982_ _3347_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__clkbuf_1
X_8721_ _4287_ vssd1 vssd1 vccd1 vccd1 _4288_ sky130_fd_sc_hd__buf_4
X_5933_ reg_data\[27\]\[23\] _2439_ _2506_ _2509_ _2512_ vssd1 vssd1 vccd1 vccd1 _2513_
+ sky130_fd_sc_hd__a2111o_1
X_5864_ reg_data\[27\]\[22\] _2439_ _2442_ _2444_ _2445_ vssd1 vssd1 vccd1 vccd1 _2446_
+ sky130_fd_sc_hd__a2111o_1
X_8652_ _3638_ _4070_ vssd1 vssd1 vccd1 vccd1 _4251_ sky130_fd_sc_hd__and2_4
X_8583_ _4214_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__clkbuf_1
X_7603_ _3206_ reg_data\[24\]\[2\] _3677_ vssd1 vssd1 vccd1 vccd1 _3680_ sky130_fd_sc_hd__mux2_1
X_4815_ reg_data\[20\]\[6\] _1312_ _1060_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__and3_1
X_5795_ reg_data\[20\]\[22\] _1918_ _1060_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__and3_1
X_7534_ reg_data\[23\]\[2\] _3133_ _3640_ vssd1 vssd1 vccd1 vccd1 _3643_ sky130_fd_sc_hd__mux2_1
X_4746_ reg_data\[26\]\[4\] _1230_ _1232_ reg_data\[29\]\[4\] vssd1 vssd1 vccd1 vccd1
+ _1364_ sky130_fd_sc_hd__a22o_1
X_4677_ reg_data\[2\]\[3\] _1002_ _1295_ _1296_ reg_data\[11\]\[3\] vssd1 vssd1 vccd1
+ vccd1 _1297_ sky130_fd_sc_hd__a32o_1
X_7465_ _3206_ reg_data\[21\]\[2\] _3603_ vssd1 vssd1 vccd1 vccd1 _3606_ sky130_fd_sc_hd__mux2_1
X_9204_ clknet_leaf_19_i_clk _0348_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6416_ reg_data\[13\]\[0\] _1177_ _1190_ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__and3_1
X_7396_ _3568_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__clkbuf_1
X_9135_ clknet_leaf_22_i_clk _0279_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6347_ _2903_ _2907_ _2909_ _2911_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__or4_1
X_6278_ reg_data\[5\]\[30\] _1085_ _2530_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__and3_1
X_9066_ clknet_leaf_44_i_clk _0210_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8017_ i_data[25] vssd1 vssd1 vccd1 vccd1 _3911_ sky130_fd_sc_hd__clkbuf_4
X_5229_ reg_data\[7\]\[12\] _1827_ _1828_ _1829_ _1830_ vssd1 vssd1 vccd1 vccd1 _1831_
+ sky130_fd_sc_hd__a2111o_1
X_8919_ clknet_leaf_25_i_clk _0063_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_9899_ clknet_leaf_73_i_clk _0969_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_4600_ reg_data\[16\]\[2\] _1219_ _1221_ reg_data\[9\]\[2\] vssd1 vssd1 vccd1 vccd1
+ _1222_ sky130_fd_sc_hd__a22o_1
X_5580_ _2170_ vssd1 vssd1 vccd1 vccd1 rdata1\[18\] sky130_fd_sc_hd__clkbuf_1
X_4531_ reg_data\[22\]\[2\] _1150_ _1152_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__and3_1
X_7250_ reg_data\[6\]\[31\] _3193_ _3455_ vssd1 vssd1 vccd1 vccd1 _3490_ sky130_fd_sc_hd__mux2_1
X_4462_ _1067_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__clkbuf_2
X_6201_ reg_data\[12\]\[28\] _2562_ _1289_ vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__and3_1
X_4393_ _1019_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__buf_2
X_7181_ _3453_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__clkbuf_1
X_6132_ _2704_ vssd1 vssd1 vccd1 vccd1 rdata1\[27\] sky130_fd_sc_hd__clkbuf_1
X_6063_ reg_data\[0\]\[26\] _2381_ _2635_ _2636_ _2637_ vssd1 vssd1 vccd1 vccd1 _2638_
+ sky130_fd_sc_hd__a2111o_1
X_5014_ _1151_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__buf_4
X_9822_ clknet_leaf_73_i_clk rdata2\[6\] vssd1 vssd1 vccd1 vccd1 r_data2\[6\] sky130_fd_sc_hd__dfxtp_2
X_6965_ _3256_ reg_data\[10\]\[26\] _3331_ vssd1 vssd1 vccd1 vccd1 _3338_ sky130_fd_sc_hd__mux2_1
X_9753_ clknet_leaf_0_i_clk _0897_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_9684_ clknet_leaf_17_i_clk _0828_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_5916_ reg_data\[3\]\[23\] _2421_ _2493_ _2494_ _2495_ vssd1 vssd1 vccd1 vccd1 _2496_
+ sky130_fd_sc_hd__a2111o_1
X_8704_ reg_data\[19\]\[24\] _3179_ _4274_ vssd1 vssd1 vccd1 vccd1 _4279_ sky130_fd_sc_hd__mux2_1
X_6896_ _3300_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__clkbuf_1
X_8635_ _4242_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__clkbuf_1
X_5847_ reg_data\[4\]\[22\] _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__and3_1
X_8566_ reg_data\[1\]\[23\] _3177_ _4202_ vssd1 vssd1 vccd1 vccd1 _4206_ sky130_fd_sc_hd__mux2_1
X_5778_ reg_data\[2\]\[21\] _1837_ _1901_ _1902_ reg_data\[11\]\[21\] vssd1 vssd1
+ vccd1 vccd1 _2362_ sky130_fd_sc_hd__a32o_1
X_7517_ _3258_ reg_data\[21\]\[27\] _3625_ vssd1 vssd1 vccd1 vccd1 _3633_ sky130_fd_sc_hd__mux2_1
X_8497_ _4169_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__clkbuf_1
X_4729_ _0999_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__clkbuf_4
X_7448_ _3595_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__clkbuf_1
X_7379_ reg_data\[3\]\[27\] _3185_ _3551_ vssd1 vssd1 vccd1 vccd1 _3559_ sky130_fd_sc_hd__mux2_1
X_9118_ clknet_leaf_3_i_clk _0262_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_9049_ clknet_leaf_13_i_clk _0193_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6750_ _3209_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__clkbuf_1
X_5701_ reg_data\[22\]\[20\] _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__and3_1
X_6681_ reg_data\[4\]\[15\] _3160_ _3150_ vssd1 vssd1 vccd1 vccd1 _3161_ sky130_fd_sc_hd__mux2_1
X_8420_ _4128_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__clkbuf_1
X_5632_ reg_data\[1\]\[19\] _1729_ _1793_ _1794_ reg_data\[15\]\[19\] vssd1 vssd1
+ vccd1 vccd1 _2221_ sky130_fd_sc_hd__a32o_1
X_5563_ reg_data\[5\]\[18\] _2097_ _1925_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__and3_1
X_8351_ _3896_ reg_data\[16\]\[18\] _4083_ vssd1 vssd1 vccd1 vccd1 _4092_ sky130_fd_sc_hd__mux2_1
X_7302_ _3518_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__clkbuf_1
X_4514_ _1093_ _1113_ _1125_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__or4_1
X_5494_ _1043_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__clkbuf_4
X_8282_ _3896_ reg_data\[15\]\[18\] _4046_ vssd1 vssd1 vccd1 vccd1 _4055_ sky130_fd_sc_hd__mux2_1
X_7233_ _3481_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__clkbuf_1
X_4445_ _1015_ _1026_ _1030_ _1033_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__and4_1
X_7164_ reg_data\[7\]\[22\] _3175_ _3442_ vssd1 vssd1 vccd1 vccd1 _3445_ sky130_fd_sc_hd__mux2_1
X_4376_ _1006_ vssd1 vssd1 vccd1 vccd1 rs2_mux\[1\] sky130_fd_sc_hd__inv_2
X_6115_ reg_data\[4\]\[27\] _2325_ _2469_ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__and3_1
X_7095_ _3248_ reg_data\[8\]\[22\] _3405_ vssd1 vssd1 vccd1 vccd1 _3408_ sky130_fd_sc_hd__mux2_1
X_6046_ reg_data\[16\]\[25\] _2449_ _2450_ reg_data\[9\]\[25\] vssd1 vssd1 vccd1 vccd1
+ _2622_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_60_i_clk clknet_3_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_9805_ clknet_leaf_50_i_clk rdata1\[21\] vssd1 vssd1 vccd1 vccd1 r_data1\[21\] sky130_fd_sc_hd__dfxtp_1
X_7997_ _3897_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_75_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_6948_ _3239_ reg_data\[10\]\[18\] _3320_ vssd1 vssd1 vccd1 vccd1 _3329_ sky130_fd_sc_hd__mux2_1
X_9736_ clknet_leaf_45_i_clk _0880_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6879_ _3291_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__clkbuf_1
X_9667_ clknet_leaf_65_i_clk _0811_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_9598_ clknet_leaf_74_i_clk _0742_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8618_ _4233_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__clkbuf_1
X_8549_ reg_data\[1\]\[15\] _3160_ _4191_ vssd1 vssd1 vccd1 vccd1 _4197_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_13_i_clk clknet_3_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_28_i_clk clknet_3_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_7920_ _3250_ reg_data\[28\]\[23\] _3844_ vssd1 vssd1 vccd1 vccd1 _3848_ sky130_fd_sc_hd__mux2_1
X_7851_ _3250_ reg_data\[27\]\[23\] _3807_ vssd1 vssd1 vccd1 vccd1 _3811_ sky130_fd_sc_hd__mux2_1
X_6802_ _3243_ reg_data\[22\]\[20\] _3244_ vssd1 vssd1 vccd1 vccd1 _3245_ sky130_fd_sc_hd__mux2_1
X_7782_ _3774_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__clkbuf_1
X_4994_ reg_data\[5\]\[9\] _1490_ _1250_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__and3_1
X_9521_ clknet_leaf_17_i_clk _0665_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6733_ _3119_ _3120_ vssd1 vssd1 vccd1 vccd1 _3196_ sky130_fd_sc_hd__nand2_1
X_6664_ i_data[10] vssd1 vssd1 vccd1 vccd1 _3149_ sky130_fd_sc_hd__buf_2
X_9452_ clknet_leaf_50_i_clk _0596_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5615_ _1034_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__clkbuf_4
X_8403_ _3879_ reg_data\[17\]\[10\] _4119_ vssd1 vssd1 vccd1 vccd1 _4120_ sky130_fd_sc_hd__mux2_1
X_6595_ _3103_ vssd1 vssd1 vccd1 vccd1 o_data2[18] sky130_fd_sc_hd__buf_2
X_9383_ clknet_leaf_56_i_clk _0527_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8334_ _4071_ vssd1 vssd1 vccd1 vccd1 _4083_ sky130_fd_sc_hd__clkbuf_4
X_5546_ reg_data\[16\]\[17\] _1843_ _1844_ reg_data\[9\]\[17\] vssd1 vssd1 vccd1 vccd1
+ _2138_ sky130_fd_sc_hd__a22o_1
X_8265_ _4034_ vssd1 vssd1 vccd1 vccd1 _4046_ sky130_fd_sc_hd__buf_4
X_5477_ reg_data\[14\]\[16\] _1693_ _1958_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__and3_1
X_4428_ rs1_mux\[2\] rs1_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__nor2_1
X_7216_ _3472_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
X_8196_ _4009_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__clkbuf_1
X_4359_ rs2\[0\] vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__inv_2
X_7147_ reg_data\[7\]\[14\] _3158_ _3431_ vssd1 vssd1 vccd1 vccd1 _3436_ sky130_fd_sc_hd__mux2_1
X_7078_ _3231_ reg_data\[8\]\[14\] _3394_ vssd1 vssd1 vccd1 vccd1 _3399_ sky130_fd_sc_hd__mux2_1
X_6029_ reg_data\[18\]\[25\] _2422_ _2120_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__and3_1
X_9719_ clknet_leaf_42_i_clk _0863_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6380_ reg_data\[25\]\[0\] _1036_ _2940_ _2941_ _2942_ vssd1 vssd1 vccd1 vccd1 _2943_
+ sky130_fd_sc_hd__a2111o_1
X_5400_ reg_data\[26\]\[15\] _1805_ _1806_ reg_data\[29\]\[15\] vssd1 vssd1 vccd1
+ vccd1 _1997_ sky130_fd_sc_hd__a22o_1
X_5331_ reg_data\[13\]\[14\] _1608_ _1257_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__and3_1
X_8050_ _3869_ reg_data\[30\]\[5\] _3926_ vssd1 vssd1 vccd1 vccd1 _3932_ sky130_fd_sc_hd__mux2_1
X_5262_ _1059_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__buf_4
X_7001_ _3357_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__clkbuf_1
X_5193_ reg_data\[27\]\[12\] _1786_ _1789_ _1792_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_
+ sky130_fd_sc_hd__a2111o_1
X_8952_ clknet_leaf_69_i_clk _0096_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8883_ clknet_leaf_15_i_clk _0027_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_7903_ _3233_ reg_data\[28\]\[15\] _3833_ vssd1 vssd1 vccd1 vccd1 _3839_ sky130_fd_sc_hd__mux2_1
X_7834_ _3233_ reg_data\[27\]\[15\] _3796_ vssd1 vssd1 vccd1 vccd1 _3802_ sky130_fd_sc_hd__mux2_1
X_7765_ _3765_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__clkbuf_1
X_6716_ _3184_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__clkbuf_1
X_4977_ reg_data\[8\]\[8\] _1214_ _1217_ reg_data\[10\]\[8\] _1586_ vssd1 vssd1 vccd1
+ vccd1 _1587_ sky130_fd_sc_hd__a221o_1
X_9504_ clknet_leaf_7_i_clk _0648_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7696_ _3231_ reg_data\[25\]\[14\] _3724_ vssd1 vssd1 vccd1 vccd1 _3729_ sky130_fd_sc_hd__mux2_1
X_9435_ clknet_leaf_71_i_clk _0579_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6647_ reg_data\[4\]\[4\] _3137_ _3129_ vssd1 vssd1 vccd1 vccd1 _3138_ sky130_fd_sc_hd__mux2_1
X_9366_ clknet_leaf_38_i_clk _0510_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6578_ r_data2\[10\] _3094_ vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__and2_1
X_5529_ reg_data\[18\]\[17\] _1816_ _2120_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__and3_1
X_8317_ _4074_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__clkbuf_1
X_9297_ clknet_leaf_35_i_clk _0441_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_8248_ _4037_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__clkbuf_1
X_8179_ _3861_ reg_data\[14\]\[1\] _3999_ vssd1 vssd1 vccd1 vccd1 _4001_ sky130_fd_sc_hd__mux2_1
X_5880_ reg_data\[21\]\[23\] _2372_ _1043_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__and3_1
X_4900_ reg_data\[25\]\[7\] _1141_ _1507_ _1508_ _1511_ vssd1 vssd1 vccd1 vccd1 _1512_
+ sky130_fd_sc_hd__a2111o_1
X_4831_ reg_data\[16\]\[6\] _1121_ _1123_ reg_data\[9\]\[6\] vssd1 vssd1 vccd1 vccd1
+ _1446_ sky130_fd_sc_hd__a22o_1
X_4762_ _1056_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__clkbuf_4
X_7550_ _3639_ vssd1 vssd1 vccd1 vccd1 _3651_ sky130_fd_sc_hd__buf_4
X_7481_ _3602_ vssd1 vssd1 vccd1 vccd1 _3614_ sky130_fd_sc_hd__buf_4
X_6501_ _3053_ vssd1 vssd1 vccd1 vccd1 o_data1[6] sky130_fd_sc_hd__buf_2
X_4693_ _1034_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__clkbuf_4
X_6432_ reg_data\[17\]\[1\] _1055_ _1040_ vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__and3_1
X_9220_ clknet_leaf_47_i_clk _0364_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_9151_ clknet_leaf_3_i_clk _0295_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8102_ _3921_ reg_data\[30\]\[30\] _3925_ vssd1 vssd1 vccd1 vccd1 _3959_ sky130_fd_sc_hd__mux2_1
X_6363_ reg_data\[13\]\[31\] _1186_ _1191_ vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__and3_1
X_6294_ _2860_ vssd1 vssd1 vccd1 vccd1 rdata1\[30\] sky130_fd_sc_hd__clkbuf_1
X_9082_ clknet_leaf_11_i_clk _0226_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_5314_ reg_data\[22\]\[14\] _1536_ _1651_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__and3_1
X_8033_ _3921_ reg_data\[9\]\[30\] _3858_ vssd1 vssd1 vccd1 vccd1 _3922_ sky130_fd_sc_hd__mux2_1
X_5245_ _1224_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__clkbuf_4
X_5176_ reg_data\[0\]\[12\] _1775_ _1776_ _1777_ _1778_ vssd1 vssd1 vccd1 vccd1 _1779_
+ sky130_fd_sc_hd__a2111o_1
X_8935_ clknet_leaf_56_i_clk _0079_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8866_ clknet_leaf_66_i_clk _0010_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8797_ _4328_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__clkbuf_1
X_7817_ _3216_ reg_data\[27\]\[7\] _3785_ vssd1 vssd1 vccd1 vccd1 _3793_ sky130_fd_sc_hd__mux2_1
X_7748_ _3756_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__clkbuf_1
X_7679_ _3214_ reg_data\[25\]\[6\] _3713_ vssd1 vssd1 vccd1 vccd1 _3720_ sky130_fd_sc_hd__mux2_1
X_9418_ clknet_leaf_53_i_clk _0562_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_9349_ clknet_leaf_58_i_clk _0493_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5030_ reg_data\[14\]\[9\] _1189_ _1193_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__and3_1
X_6981_ reg_data\[0\]\[1\] _3131_ _3345_ vssd1 vssd1 vccd1 vccd1 _3347_ sky130_fd_sc_hd__mux2_1
X_5932_ reg_data\[1\]\[23\] _2510_ _2511_ reg_data\[15\]\[23\] vssd1 vssd1 vccd1 vccd1
+ _2512_ sky130_fd_sc_hd__a22o_1
X_8720_ _3491_ _3820_ vssd1 vssd1 vccd1 vccd1 _4287_ sky130_fd_sc_hd__or2_4
X_8651_ _4250_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__clkbuf_1
X_5863_ reg_data\[1\]\[22\] _1904_ _1905_ reg_data\[15\]\[22\] vssd1 vssd1 vccd1 vccd1
+ _2445_ sky130_fd_sc_hd__a22o_1
X_5794_ reg_data\[18\]\[22\] _2261_ _2090_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__and3_1
X_8582_ reg_data\[1\]\[31\] _3193_ _4179_ vssd1 vssd1 vccd1 vccd1 _4214_ sky130_fd_sc_hd__mux2_1
X_7602_ _3679_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__clkbuf_1
X_4814_ reg_data\[18\]\[6\] _1055_ _1064_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__and3_1
X_4745_ reg_data\[8\]\[4\] _1214_ _1217_ reg_data\[10\]\[4\] _1362_ vssd1 vssd1 vccd1
+ vccd1 _1363_ sky130_fd_sc_hd__a221o_1
X_7533_ _3642_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__clkbuf_1
X_4676_ _1200_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__buf_4
X_7464_ _3605_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__clkbuf_1
X_9203_ clknet_leaf_18_i_clk _0347_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6415_ reg_data\[0\]\[0\] _1173_ _2974_ _2975_ _2976_ vssd1 vssd1 vccd1 vccd1 _2977_
+ sky130_fd_sc_hd__a2111o_1
X_7395_ _3206_ reg_data\[20\]\[2\] _3565_ vssd1 vssd1 vccd1 vccd1 _3568_ sky130_fd_sc_hd__mux2_1
X_9134_ clknet_leaf_29_i_clk _0278_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6346_ reg_data\[24\]\[31\] _2409_ _2410_ reg_data\[28\]\[31\] _2910_ vssd1 vssd1
+ vccd1 vccd1 _2911_ sky130_fd_sc_hd__a221o_1
X_9065_ clknet_leaf_44_i_clk _0209_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_8016_ _3910_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__clkbuf_1
X_6277_ reg_data\[4\]\[30\] _2325_ _2469_ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__and3_1
X_5228_ reg_data\[12\]\[12\] _1354_ _1226_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__and3_1
X_5159_ _1754_ _1758_ _1760_ _1762_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__or4_1
X_8918_ clknet_leaf_24_i_clk _0062_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_9898_ clknet_leaf_75_i_clk _0968_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8849_ _4355_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__clkbuf_1
X_4530_ _1151_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__clkbuf_4
X_4461_ reg_data\[12\]\[2\] _1082_ _1083_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__and3_1
X_6200_ reg_data\[14\]\[28\] _2301_ _1344_ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__and3_1
X_7180_ reg_data\[7\]\[30\] _3191_ _3419_ vssd1 vssd1 vccd1 vccd1 _3453_ sky130_fd_sc_hd__mux2_1
X_6131_ _2695_ _2699_ _2701_ _2703_ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__or4_1
X_4392_ _0995_ i_rs1[4] _1016_ _1018_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__o31a_1
X_6062_ reg_data\[5\]\[26\] _2097_ _2530_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__and3_1
X_5013_ _1621_ vssd1 vssd1 vccd1 vccd1 rdata1\[9\] sky130_fd_sc_hd__clkbuf_1
X_9821_ clknet_leaf_62_i_clk rdata2\[5\] vssd1 vssd1 vccd1 vccd1 r_data2\[5\] sky130_fd_sc_hd__dfxtp_1
X_6964_ _3337_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__clkbuf_1
X_9752_ clknet_leaf_69_i_clk _0896_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_9683_ clknet_leaf_17_i_clk _0827_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5915_ reg_data\[20\]\[23\] _2234_ _1743_ vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__and3_1
X_6895_ reg_data\[2\]\[26\] _3183_ _3293_ vssd1 vssd1 vccd1 vccd1 _3300_ sky130_fd_sc_hd__mux2_1
X_8703_ _4278_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__clkbuf_1
X_8634_ _3907_ reg_data\[12\]\[23\] _4238_ vssd1 vssd1 vccd1 vccd1 _4242_ sky130_fd_sc_hd__mux2_1
X_5846_ reg_data\[6\]\[22\] _1951_ _2237_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__and3_1
X_8565_ _4205_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__clkbuf_1
X_5777_ reg_data\[23\]\[21\] _1834_ _1835_ reg_data\[19\]\[21\] vssd1 vssd1 vccd1
+ vccd1 _2361_ sky130_fd_sc_hd__a22o_1
X_7516_ _3632_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__clkbuf_1
X_8496_ _3905_ reg_data\[18\]\[22\] _4166_ vssd1 vssd1 vccd1 vccd1 _4169_ sky130_fd_sc_hd__mux2_1
X_4728_ reg_data\[3\]\[4\] _1158_ _1341_ _1343_ _1345_ vssd1 vssd1 vccd1 vccd1 _1346_
+ sky130_fd_sc_hd__a2111o_1
X_7447_ _3258_ reg_data\[20\]\[27\] _3587_ vssd1 vssd1 vccd1 vccd1 _3595_ sky130_fd_sc_hd__mux2_1
X_4659_ reg_data\[30\]\[3\] _1162_ _1164_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__and3_1
X_7378_ _3558_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__clkbuf_1
X_6329_ reg_data\[3\]\[31\] _2376_ _2891_ _2892_ _2893_ vssd1 vssd1 vccd1 vccd1 _2894_
+ sky130_fd_sc_hd__a2111o_1
X_9117_ clknet_leaf_3_i_clk _0261_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_9048_ clknet_leaf_13_i_clk _0192_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_5__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5700_ _1151_ vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__buf_2
X_6680_ i_data[15] vssd1 vssd1 vccd1 vccd1 _3160_ sky130_fd_sc_hd__clkbuf_4
X_5631_ reg_data\[2\]\[19\] _2219_ _1790_ _1791_ reg_data\[11\]\[19\] vssd1 vssd1
+ vccd1 vccd1 _2220_ sky130_fd_sc_hd__a32o_1
X_5562_ reg_data\[4\]\[18\] _1718_ _1863_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__and3_1
X_8350_ _4091_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__clkbuf_1
X_7301_ reg_data\[5\]\[22\] _3175_ _3515_ vssd1 vssd1 vccd1 vccd1 _3518_ sky130_fd_sc_hd__mux2_1
X_8281_ _4054_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__clkbuf_1
X_4513_ reg_data\[24\]\[2\] _1127_ _1130_ reg_data\[28\]\[2\] _1135_ vssd1 vssd1 vccd1
+ vccd1 _1136_ sky130_fd_sc_hd__a221o_1
X_7232_ reg_data\[6\]\[22\] _3175_ _3478_ vssd1 vssd1 vccd1 vccd1 _3481_ sky130_fd_sc_hd__mux2_1
X_5493_ _1034_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__clkbuf_4
X_4444_ _1019_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__buf_2
X_7163_ _3444_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__clkbuf_1
X_4375_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__buf_2
X_6114_ reg_data\[6\]\[27\] _2207_ _2323_ vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__and3_1
X_7094_ _3407_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__clkbuf_1
X_6045_ reg_data\[27\]\[25\] _2439_ _2618_ _2619_ _2620_ vssd1 vssd1 vccd1 vccd1 _2621_
+ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_9_i_clk clknet_3_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_9804_ clknet_leaf_50_i_clk rdata1\[20\] vssd1 vssd1 vccd1 vccd1 r_data1\[20\] sky130_fd_sc_hd__dfxtp_1
X_7996_ _3896_ reg_data\[9\]\[18\] _3880_ vssd1 vssd1 vccd1 vccd1 _3897_ sky130_fd_sc_hd__mux2_1
X_9735_ clknet_leaf_8_i_clk _0879_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6947_ _3328_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__clkbuf_1
X_6878_ reg_data\[2\]\[18\] _3166_ _3282_ vssd1 vssd1 vccd1 vccd1 _3291_ sky130_fd_sc_hd__mux2_1
X_9666_ clknet_leaf_65_i_clk _0810_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_5829_ _1133_ vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__clkbuf_4
X_9597_ clknet_leaf_70_i_clk _0741_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_8617_ _3890_ reg_data\[12\]\[15\] _4227_ vssd1 vssd1 vccd1 vccd1 _4233_ sky130_fd_sc_hd__mux2_1
X_8548_ _4196_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__clkbuf_1
X_8479_ _3888_ reg_data\[18\]\[14\] _4155_ vssd1 vssd1 vccd1 vccd1 _4160_ sky130_fd_sc_hd__mux2_1
X_7850_ _3810_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__clkbuf_1
X_6801_ _3201_ vssd1 vssd1 vccd1 vccd1 _3244_ sky130_fd_sc_hd__buf_4
X_7781_ _3248_ reg_data\[26\]\[22\] _3771_ vssd1 vssd1 vccd1 vccd1 _3774_ sky130_fd_sc_hd__mux2_1
X_4993_ reg_data\[4\]\[9\] _1074_ _1248_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__and3_1
X_9520_ clknet_leaf_18_i_clk _0664_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6732_ i_data[0] vssd1 vssd1 vccd1 vccd1 _3195_ sky130_fd_sc_hd__clkbuf_4
X_9451_ clknet_leaf_63_i_clk _0595_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6663_ _3148_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__clkbuf_1
X_5614_ reg_data\[20\]\[19\] _1918_ _1060_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__and3_1
X_8402_ _4107_ vssd1 vssd1 vccd1 vccd1 _4119_ sky130_fd_sc_hd__buf_6
X_9382_ clknet_leaf_54_i_clk _0526_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6594_ r_data2\[18\] _3094_ vssd1 vssd1 vccd1 vccd1 _3103_ sky130_fd_sc_hd__and2_1
X_5545_ reg_data\[27\]\[17\] _1833_ _2134_ _2135_ _2136_ vssd1 vssd1 vccd1 vccd1 _2137_
+ sky130_fd_sc_hd__a2111o_1
X_8333_ _4082_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__clkbuf_1
X_8264_ _4045_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__clkbuf_1
X_5476_ reg_data\[13\]\[16\] _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__and3_1
X_7215_ reg_data\[6\]\[14\] _3158_ _3467_ vssd1 vssd1 vccd1 vccd1 _3472_ sky130_fd_sc_hd__mux2_1
X_8195_ _3877_ reg_data\[14\]\[9\] _3999_ vssd1 vssd1 vccd1 vccd1 _4009_ sky130_fd_sc_hd__mux2_1
X_4427_ reg_data\[25\]\[2\] _1037_ _1041_ _1045_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_
+ sky130_fd_sc_hd__a2111o_1
X_7146_ _3435_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_1
X_7077_ _3398_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
X_6028_ reg_data\[25\]\[25\] _2416_ _2601_ _2602_ _2603_ vssd1 vssd1 vccd1 vccd1 _2604_
+ sky130_fd_sc_hd__a2111o_1
X_7979_ _3885_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__clkbuf_1
X_9718_ clknet_leaf_39_i_clk _0862_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_9649_ clknet_leaf_21_i_clk _0793_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_5330_ reg_data\[12\]\[14\] _1381_ _1606_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__and3_1
X_5261_ reg_data\[6\]\[13\] _1600_ _1716_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__and3_1
X_7000_ reg_data\[0\]\[10\] _3149_ _3356_ vssd1 vssd1 vccd1 vccd1 _3357_ sky130_fd_sc_hd__mux2_1
X_5192_ reg_data\[1\]\[12\] _1729_ _1793_ _1794_ reg_data\[15\]\[12\] vssd1 vssd1
+ vccd1 vccd1 _1795_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_74_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_8951_ clknet_leaf_41_i_clk _0095_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_7902_ _3838_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__clkbuf_1
X_8882_ clknet_leaf_20_i_clk _0026_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_7833_ _3801_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_12_i_clk clknet_3_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_7764_ _3231_ reg_data\[26\]\[14\] _3760_ vssd1 vssd1 vccd1 vccd1 _3765_ sky130_fd_sc_hd__mux2_1
X_6715_ reg_data\[4\]\[26\] _3183_ _3171_ vssd1 vssd1 vccd1 vccd1 _3184_ sky130_fd_sc_hd__mux2_1
X_4976_ reg_data\[16\]\[8\] _1219_ _1221_ reg_data\[9\]\[8\] vssd1 vssd1 vccd1 vccd1
+ _1586_ sky130_fd_sc_hd__a22o_1
X_9503_ clknet_leaf_4_i_clk _0647_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_7695_ _3728_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__clkbuf_1
X_9434_ clknet_leaf_70_i_clk _0578_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6646_ i_data[4] vssd1 vssd1 vccd1 vccd1 _3137_ sky130_fd_sc_hd__clkbuf_4
X_9365_ clknet_leaf_34_i_clk _0509_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_27_i_clk clknet_3_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_6577_ _3082_ vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__dlymetal6s2s_1
X_5528_ _1167_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__clkbuf_4
X_8316_ _3861_ reg_data\[16\]\[1\] _4072_ vssd1 vssd1 vccd1 vccd1 _4074_ sky130_fd_sc_hd__mux2_1
X_9296_ clknet_leaf_34_i_clk _0440_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_8247_ _3861_ reg_data\[15\]\[1\] _4035_ vssd1 vssd1 vccd1 vccd1 _4037_ sky130_fd_sc_hd__mux2_1
X_5459_ reg_data\[24\]\[16\] _1803_ _1804_ reg_data\[28\]\[16\] _2053_ vssd1 vssd1
+ vccd1 vccd1 _2054_ sky130_fd_sc_hd__a221o_1
X_8178_ _4000_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__clkbuf_1
X_7129_ _3426_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__clkbuf_1
X_4830_ reg_data\[27\]\[6\] _1096_ _1442_ _1443_ _1444_ vssd1 vssd1 vccd1 vccd1 _1445_
+ sky130_fd_sc_hd__a2111o_1
X_4761_ reg_data\[0\]\[5\] _1070_ _1375_ _1376_ _1377_ vssd1 vssd1 vccd1 vccd1 _1378_
+ sky130_fd_sc_hd__a2111o_1
X_6500_ r_data1\[6\] _3046_ vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__and2_1
X_7480_ _3613_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__clkbuf_1
X_4692_ reg_data\[18\]\[4\] _1055_ _1064_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__and3_1
X_6431_ reg_data\[22\]\[1\] _1097_ _1047_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__and3_1
X_6362_ reg_data\[14\]\[31\] _1177_ _1164_ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__and3_1
X_9150_ clknet_leaf_3_i_clk _0294_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8101_ _3958_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__clkbuf_1
X_5313_ _1912_ vssd1 vssd1 vccd1 vccd1 rdata2\[13\] sky130_fd_sc_hd__clkbuf_1
X_6293_ _2851_ _2855_ _2857_ _2859_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__or4_1
X_9081_ clknet_leaf_12_i_clk _0225_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8032_ i_data[30] vssd1 vssd1 vccd1 vccd1 _3921_ sky130_fd_sc_hd__buf_4
X_5244_ reg_data\[8\]\[12\] _1841_ _1842_ reg_data\[10\]\[12\] _1845_ vssd1 vssd1
+ vccd1 vccd1 _1846_ sky130_fd_sc_hd__a221o_1
X_5175_ reg_data\[5\]\[12\] _1490_ _1250_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__and3_1
X_8934_ clknet_leaf_56_i_clk _0078_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8865_ clknet_leaf_2_i_clk _0009_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_7816_ _3792_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__clkbuf_1
X_8796_ reg_data\[11\]\[3\] i_data[3] _4324_ vssd1 vssd1 vccd1 vccd1 _4328_ sky130_fd_sc_hd__mux2_1
X_7747_ _3214_ reg_data\[26\]\[6\] _3749_ vssd1 vssd1 vccd1 vccd1 _3756_ sky130_fd_sc_hd__mux2_1
X_4959_ reg_data\[20\]\[8\] _1166_ _1180_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__and3_1
X_7678_ _3719_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__clkbuf_1
X_9417_ clknet_leaf_58_i_clk _0561_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6629_ _3122_ _3123_ vssd1 vssd1 vccd1 vccd1 _3124_ sky130_fd_sc_hd__nand2_1
X_9348_ clknet_leaf_59_i_clk _0492_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_9279_ clknet_leaf_72_i_clk _0423_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6980_ _3346_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__clkbuf_1
X_5931_ _1203_ vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__buf_4
X_8650_ _3923_ reg_data\[12\]\[31\] _4215_ vssd1 vssd1 vccd1 vccd1 _4250_ sky130_fd_sc_hd__mux2_1
X_5862_ reg_data\[2\]\[22\] _2443_ _1901_ _1902_ reg_data\[11\]\[22\] vssd1 vssd1
+ vccd1 vccd1 _2444_ sky130_fd_sc_hd__a32o_1
X_5793_ _1053_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__clkbuf_4
X_8581_ _4213_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__clkbuf_1
X_7601_ _3204_ reg_data\[24\]\[1\] _3677_ vssd1 vssd1 vccd1 vccd1 _3679_ sky130_fd_sc_hd__mux2_1
X_4813_ reg_data\[25\]\[6\] _1037_ _1425_ _1426_ _1427_ vssd1 vssd1 vccd1 vccd1 _1428_
+ sky130_fd_sc_hd__a2111o_1
X_4744_ reg_data\[16\]\[4\] _1219_ _1221_ reg_data\[9\]\[4\] vssd1 vssd1 vccd1 vccd1
+ _1362_ sky130_fd_sc_hd__a22o_1
X_7532_ reg_data\[23\]\[1\] _3131_ _3640_ vssd1 vssd1 vccd1 vccd1 _3642_ sky130_fd_sc_hd__mux2_1
X_9202_ clknet_leaf_30_i_clk _0346_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_4675_ _1168_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__buf_4
X_7463_ _3204_ reg_data\[21\]\[1\] _3603_ vssd1 vssd1 vccd1 vccd1 _3605_ sky130_fd_sc_hd__mux2_1
X_6414_ reg_data\[5\]\[0\] _1189_ _1338_ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__and3_1
X_7394_ _3567_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__clkbuf_1
X_6345_ reg_data\[26\]\[31\] _2411_ _2412_ reg_data\[29\]\[31\] vssd1 vssd1 vccd1
+ vccd1 _2910_ sky130_fd_sc_hd__a22o_1
X_9133_ clknet_leaf_27_i_clk _0277_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6276_ reg_data\[6\]\[30\] _1020_ _2323_ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__and3_1
X_9064_ clknet_leaf_46_i_clk _0208_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_8015_ _3909_ reg_data\[9\]\[24\] _3901_ vssd1 vssd1 vccd1 vccd1 _3910_ sky130_fd_sc_hd__mux2_1
X_5227_ reg_data\[14\]\[12\] _1693_ _1193_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__and3_1
X_5158_ reg_data\[24\]\[11\] _1225_ _1228_ reg_data\[28\]\[11\] _1761_ vssd1 vssd1
+ vccd1 vccd1 _1762_ sky130_fd_sc_hd__a221o_1
X_5089_ reg_data\[14\]\[10\] _1354_ _1193_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__and3_1
X_8917_ clknet_leaf_21_i_clk _0061_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_9897_ clknet_leaf_77_i_clk _0967_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8848_ reg_data\[11\]\[28\] i_data[28] _4346_ vssd1 vssd1 vccd1 vccd1 _4355_ sky130_fd_sc_hd__mux2_1
X_8779_ _4318_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__clkbuf_1
X_4460_ _1015_ _1026_ rs1_mux\[2\] rs1_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__and4_2
X_4391_ _0995_ _1016_ _1017_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__o21ai_1
X_6130_ reg_data\[24\]\[27\] _2409_ _2410_ reg_data\[28\]\[27\] _2702_ vssd1 vssd1
+ vccd1 vccd1 _2703_ sky130_fd_sc_hd__a221o_1
X_6061_ reg_data\[4\]\[26\] _2325_ _2469_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__and3_1
X_5012_ _1611_ _1616_ _1618_ _1620_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__or4_1
X_9820_ clknet_leaf_59_i_clk rdata2\[4\] vssd1 vssd1 vccd1 vccd1 r_data2\[4\] sky130_fd_sc_hd__dfxtp_1
X_6963_ _3254_ reg_data\[10\]\[25\] _3331_ vssd1 vssd1 vccd1 vccd1 _3337_ sky130_fd_sc_hd__mux2_1
X_9751_ clknet_leaf_13_i_clk _0895_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_9682_ clknet_leaf_18_i_clk _0826_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_5914_ reg_data\[30\]\[23\] _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__and3_1
X_6894_ _3299_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__clkbuf_1
X_8702_ reg_data\[19\]\[23\] _3177_ _4274_ vssd1 vssd1 vccd1 vccd1 _4278_ sky130_fd_sc_hd__mux2_1
X_8633_ _4241_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__clkbuf_1
X_5845_ _1173_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__clkbuf_4
X_5776_ _2347_ _2351_ _2355_ _2359_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__or4_2
X_8564_ reg_data\[1\]\[22\] _3175_ _4202_ vssd1 vssd1 vccd1 vccd1 _4205_ sky130_fd_sc_hd__mux2_1
X_7515_ _3256_ reg_data\[21\]\[26\] _3625_ vssd1 vssd1 vccd1 vccd1 _3632_ sky130_fd_sc_hd__mux2_1
X_8495_ _4168_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__clkbuf_1
X_4727_ reg_data\[30\]\[4\] _1166_ _1344_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__and3_1
X_7446_ _3594_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__clkbuf_1
X_4658_ reg_data\[18\]\[3\] _1159_ _1168_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__and3_1
X_7377_ reg_data\[3\]\[26\] _3183_ _3551_ vssd1 vssd1 vccd1 vccd1 _3558_ sky130_fd_sc_hd__mux2_1
X_4589_ reg_data\[27\]\[2\] _1199_ _1201_ _1204_ _1210_ vssd1 vssd1 vccd1 vccd1 _1211_
+ sky130_fd_sc_hd__a2111o_1
X_9116_ clknet_leaf_4_i_clk _0260_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6328_ reg_data\[20\]\[31\] _1046_ _2035_ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__and3_1
X_6259_ reg_data\[2\]\[29\] _2443_ _2507_ _2508_ reg_data\[11\]\[29\] vssd1 vssd1
+ vccd1 vccd1 _2827_ sky130_fd_sc_hd__a32o_1
X_9047_ clknet_leaf_43_i_clk _0191_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5630_ _1089_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__buf_4
X_5561_ reg_data\[6\]\[18\] _1600_ _1716_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__and3_1
X_7300_ _3517_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__clkbuf_1
X_5492_ reg_data\[17\]\[17\] _1766_ _1708_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__and3_1
X_8280_ _3894_ reg_data\[15\]\[17\] _4046_ vssd1 vssd1 vccd1 vccd1 _4054_ sky130_fd_sc_hd__mux2_1
X_4512_ reg_data\[26\]\[2\] _1132_ _1134_ reg_data\[29\]\[2\] vssd1 vssd1 vccd1 vccd1
+ _1135_ sky130_fd_sc_hd__a22o_1
X_7231_ _3480_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__clkbuf_1
X_4443_ reg_data\[3\]\[2\] _1054_ _1057_ _1061_ _1065_ vssd1 vssd1 vccd1 vccd1 _1066_
+ sky130_fd_sc_hd__a2111o_1
X_4374_ _0994_ rs2\[1\] _1003_ _1004_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__a2bb2o_1
X_7162_ reg_data\[7\]\[21\] _3173_ _3442_ vssd1 vssd1 vccd1 vccd1 _3444_ sky130_fd_sc_hd__mux2_1
X_6113_ reg_data\[3\]\[27\] _2376_ _2683_ _2684_ _2685_ vssd1 vssd1 vccd1 vccd1 _2686_
+ sky130_fd_sc_hd__a2111o_1
X_7093_ _3246_ reg_data\[8\]\[21\] _3405_ vssd1 vssd1 vccd1 vccd1 _3407_ sky130_fd_sc_hd__mux2_1
X_6044_ reg_data\[1\]\[25\] _2510_ _2511_ reg_data\[15\]\[25\] vssd1 vssd1 vccd1 vccd1
+ _2620_ sky130_fd_sc_hd__a22o_1
X_7995_ i_data[18] vssd1 vssd1 vccd1 vccd1 _3896_ sky130_fd_sc_hd__clkbuf_4
X_9803_ clknet_leaf_58_i_clk rdata1\[19\] vssd1 vssd1 vccd1 vccd1 r_data1\[19\] sky130_fd_sc_hd__dfxtp_1
X_6946_ _3237_ reg_data\[10\]\[17\] _3320_ vssd1 vssd1 vccd1 vccd1 _3328_ sky130_fd_sc_hd__mux2_1
X_9734_ clknet_leaf_65_i_clk _0878_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6877_ _3290_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__clkbuf_1
X_9665_ clknet_leaf_5_i_clk _0809_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5828_ _1131_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__clkbuf_4
X_9596_ clknet_leaf_74_i_clk _0740_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_8616_ _4232_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__clkbuf_1
X_8547_ reg_data\[1\]\[14\] _3158_ _4191_ vssd1 vssd1 vccd1 vccd1 _4196_ sky130_fd_sc_hd__mux2_1
X_5759_ _2343_ vssd1 vssd1 vccd1 vccd1 rdata1\[21\] sky130_fd_sc_hd__clkbuf_1
X_8478_ _4159_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__clkbuf_1
X_7429_ _3585_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__clkbuf_1
X_6800_ i_data[20] vssd1 vssd1 vccd1 vccd1 _3243_ sky130_fd_sc_hd__clkbuf_4
X_4992_ reg_data\[6\]\[9\] _1600_ _1048_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__and3_1
X_7780_ _3773_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__clkbuf_1
X_6731_ _3194_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__clkbuf_1
X_6662_ reg_data\[4\]\[9\] _3147_ _3129_ vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__mux2_1
X_9450_ clknet_leaf_51_i_clk _0594_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_5613_ reg_data\[18\]\[19\] _1656_ _2090_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__and3_1
X_9381_ clknet_leaf_58_i_clk _0525_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8401_ _4118_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__clkbuf_1
X_6593_ _3102_ vssd1 vssd1 vccd1 vccd1 o_data2[17] sky130_fd_sc_hd__buf_2
X_8332_ _3877_ reg_data\[16\]\[9\] _4072_ vssd1 vssd1 vccd1 vccd1 _4082_ sky130_fd_sc_hd__mux2_1
X_5544_ reg_data\[1\]\[17\] _1904_ _1905_ reg_data\[15\]\[17\] vssd1 vssd1 vccd1 vccd1
+ _2136_ sky130_fd_sc_hd__a22o_1
X_8263_ _3877_ reg_data\[15\]\[9\] _4035_ vssd1 vssd1 vccd1 vccd1 _4045_ sky130_fd_sc_hd__mux2_1
X_5475_ reg_data\[0\]\[16\] _1821_ _2064_ _2067_ _2068_ vssd1 vssd1 vccd1 vccd1 _2069_
+ sky130_fd_sc_hd__a2111o_1
X_7214_ _3471_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
X_8194_ _4008_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__clkbuf_1
X_4426_ reg_data\[22\]\[2\] _1046_ _1048_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__and3_1
X_7145_ reg_data\[7\]\[13\] _3156_ _3431_ vssd1 vssd1 vccd1 vccd1 _3435_ sky130_fd_sc_hd__mux2_1
X_7076_ _3229_ reg_data\[8\]\[13\] _3394_ vssd1 vssd1 vccd1 vccd1 _3398_ sky130_fd_sc_hd__mux2_1
X_6027_ reg_data\[17\]\[25\] _2117_ _1148_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__and3_1
X_7978_ _3884_ reg_data\[9\]\[12\] _3880_ vssd1 vssd1 vccd1 vccd1 _3885_ sky130_fd_sc_hd__mux2_1
X_9717_ clknet_leaf_36_i_clk _0861_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6929_ _3220_ reg_data\[10\]\[9\] _3309_ vssd1 vssd1 vccd1 vccd1 _3319_ sky130_fd_sc_hd__mux2_1
X_9648_ clknet_leaf_22_i_clk _0792_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_9579_ clknet_leaf_59_i_clk _0723_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_8_i_clk clknet_3_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5260_ reg_data\[3\]\[13\] _1770_ _1858_ _1859_ _1860_ vssd1 vssd1 vccd1 vccd1 _1861_
+ sky130_fd_sc_hd__a2111o_1
X_5191_ _1110_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__buf_4
X_8950_ clknet_leaf_39_i_clk _0094_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_7901_ _3231_ reg_data\[28\]\[14\] _3833_ vssd1 vssd1 vccd1 vccd1 _3838_ sky130_fd_sc_hd__mux2_1
X_8881_ clknet_leaf_23_i_clk _0025_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_7832_ _3231_ reg_data\[27\]\[14\] _3796_ vssd1 vssd1 vccd1 vccd1 _3801_ sky130_fd_sc_hd__mux2_1
X_4975_ reg_data\[27\]\[8\] _1199_ _1582_ _1583_ _1584_ vssd1 vssd1 vccd1 vccd1 _1585_
+ sky130_fd_sc_hd__a2111o_1
X_7763_ _3764_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__clkbuf_1
X_6714_ i_data[26] vssd1 vssd1 vccd1 vccd1 _3183_ sky130_fd_sc_hd__buf_4
X_9502_ clknet_leaf_4_i_clk _0646_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_9433_ clknet_leaf_67_i_clk _0577_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_7694_ _3229_ reg_data\[25\]\[13\] _3724_ vssd1 vssd1 vccd1 vccd1 _3728_ sky130_fd_sc_hd__mux2_1
X_6645_ _3136_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__clkbuf_1
X_9364_ clknet_leaf_31_i_clk _0508_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6576_ _3093_ vssd1 vssd1 vccd1 vccd1 o_data2[9] sky130_fd_sc_hd__buf_2
X_9295_ clknet_leaf_33_i_clk _0439_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_5527_ reg_data\[25\]\[17\] _1810_ _2115_ _2116_ _2118_ vssd1 vssd1 vccd1 vccd1 _2119_
+ sky130_fd_sc_hd__a2111o_1
X_8315_ _4073_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__clkbuf_1
X_8246_ _4036_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__clkbuf_1
X_5458_ reg_data\[26\]\[16\] _1805_ _1806_ reg_data\[29\]\[16\] vssd1 vssd1 vccd1
+ vccd1 _2053_ sky130_fd_sc_hd__a22o_1
X_4409_ _0994_ _1016_ _1031_ _1032_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__a31o_2
X_8177_ _3857_ reg_data\[14\]\[0\] _3999_ vssd1 vssd1 vccd1 vccd1 _4000_ sky130_fd_sc_hd__mux2_1
X_5389_ _1067_ vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__clkbuf_4
X_7128_ reg_data\[7\]\[5\] _3139_ _3420_ vssd1 vssd1 vccd1 vccd1 _3426_ sky130_fd_sc_hd__mux2_1
X_7059_ _3212_ reg_data\[8\]\[5\] _3383_ vssd1 vssd1 vccd1 vccd1 _3389_ sky130_fd_sc_hd__mux2_1
X_4760_ reg_data\[5\]\[5\] _1076_ _1250_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__and3_1
X_4691_ reg_data\[25\]\[4\] _1037_ _1307_ _1308_ _1309_ vssd1 vssd1 vccd1 vccd1 _1310_
+ sky130_fd_sc_hd__a2111o_1
X_6430_ _2991_ vssd1 vssd1 vccd1 vccd1 rdata2\[0\] sky130_fd_sc_hd__clkbuf_1
X_6361_ reg_data\[0\]\[31\] _2427_ _2922_ _2923_ _2924_ vssd1 vssd1 vccd1 vccd1 _2925_
+ sky130_fd_sc_hd__a2111o_1
X_8100_ _3919_ reg_data\[30\]\[29\] _3948_ vssd1 vssd1 vccd1 vccd1 _3958_ sky130_fd_sc_hd__mux2_1
X_5312_ _1899_ _1907_ _1909_ _1911_ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__or4_1
X_6292_ reg_data\[24\]\[30\] _2409_ _2410_ reg_data\[28\]\[30\] _2858_ vssd1 vssd1
+ vccd1 vccd1 _2859_ sky130_fd_sc_hd__a221o_1
X_9080_ clknet_leaf_13_i_clk _0224_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8031_ _3920_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__clkbuf_1
X_5243_ reg_data\[16\]\[12\] _1843_ _1844_ reg_data\[9\]\[12\] vssd1 vssd1 vccd1 vccd1
+ _1845_ sky130_fd_sc_hd__a22o_1
X_5174_ reg_data\[4\]\[12\] _1718_ _1248_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__and3_1
X_8933_ clknet_leaf_57_i_clk _0077_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8864_ clknet_leaf_2_i_clk _0008_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7815_ _3214_ reg_data\[27\]\[6\] _3785_ vssd1 vssd1 vccd1 vccd1 _3792_ sky130_fd_sc_hd__mux2_1
X_8795_ _4327_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__clkbuf_1
X_7746_ _3755_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__clkbuf_1
X_4958_ reg_data\[30\]\[8\] _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__and3_1
X_4889_ reg_data\[16\]\[7\] _1121_ _1123_ reg_data\[9\]\[7\] vssd1 vssd1 vccd1 vccd1
+ _1502_ sky130_fd_sc_hd__a22o_1
X_7677_ _3212_ reg_data\[25\]\[5\] _3713_ vssd1 vssd1 vccd1 vccd1 _3719_ sky130_fd_sc_hd__mux2_1
X_9416_ clknet_leaf_53_i_clk _0560_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6628_ i_rd[3] _3119_ vssd1 vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__nand2_1
X_9347_ clknet_leaf_60_i_clk _0491_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6559_ r_data2\[1\] _3083_ vssd1 vssd1 vccd1 vccd1 _3085_ sky130_fd_sc_hd__and2_1
X_9278_ clknet_leaf_72_i_clk _0422_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8229_ _3911_ reg_data\[14\]\[25\] _4021_ vssd1 vssd1 vccd1 vccd1 _4027_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_73_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_11_i_clk clknet_3_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_26_i_clk clknet_3_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5930_ _1202_ vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__buf_4
X_5861_ _1001_ vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__clkbuf_4
X_7600_ _3678_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__clkbuf_1
X_5792_ reg_data\[25\]\[22\] _2370_ _2371_ _2373_ _2374_ vssd1 vssd1 vccd1 vccd1 _2375_
+ sky130_fd_sc_hd__a2111o_1
X_8580_ reg_data\[1\]\[30\] _3191_ _4179_ vssd1 vssd1 vccd1 vccd1 _4213_ sky130_fd_sc_hd__mux2_1
X_4812_ reg_data\[21\]\[6\] _1046_ _1240_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__and3_1
X_4743_ reg_data\[27\]\[4\] _1199_ _1358_ _1359_ _1360_ vssd1 vssd1 vccd1 vccd1 _1361_
+ sky130_fd_sc_hd__a2111o_1
X_7531_ _3641_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__clkbuf_1
X_7462_ _3604_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__clkbuf_1
X_9201_ clknet_leaf_21_i_clk _0345_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6413_ reg_data\[4\]\[0\] _1175_ _1342_ vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__and3_1
X_4674_ reg_data\[23\]\[3\] _1206_ _1209_ reg_data\[19\]\[3\] vssd1 vssd1 vccd1 vccd1
+ _1294_ sky130_fd_sc_hd__a22o_1
X_7393_ _3204_ reg_data\[20\]\[1\] _3565_ vssd1 vssd1 vccd1 vccd1 _3567_ sky130_fd_sc_hd__mux2_1
X_6344_ reg_data\[8\]\[31\] _2403_ _2404_ reg_data\[10\]\[31\] _2908_ vssd1 vssd1
+ vccd1 vccd1 _2909_ sky130_fd_sc_hd__a221o_1
X_9132_ clknet_leaf_27_i_clk _0276_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6275_ reg_data\[3\]\[30\] _2376_ _2839_ _2840_ _2841_ vssd1 vssd1 vccd1 vccd1 _2842_
+ sky130_fd_sc_hd__a2111o_1
X_9063_ clknet_leaf_46_i_clk _0207_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8014_ i_data[24] vssd1 vssd1 vccd1 vccd1 _3909_ sky130_fd_sc_hd__clkbuf_4
X_5226_ reg_data\[13\]\[12\] _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__and3_1
X_5157_ reg_data\[26\]\[11\] _1230_ _1232_ reg_data\[29\]\[11\] vssd1 vssd1 vccd1
+ vccd1 _1761_ sky130_fd_sc_hd__a22o_1
X_5088_ reg_data\[12\]\[10\] _1693_ _1289_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__and3_1
X_8916_ clknet_leaf_21_i_clk _0060_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_9896_ clknet_leaf_75_i_clk _0966_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8847_ _4354_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__clkbuf_1
X_8778_ _3915_ reg_data\[29\]\[27\] _4310_ vssd1 vssd1 vccd1 vccd1 _4318_ sky130_fd_sc_hd__mux2_1
X_7729_ _3264_ reg_data\[25\]\[30\] _3712_ vssd1 vssd1 vccd1 vccd1 _3746_ sky130_fd_sc_hd__mux2_1
X_4390_ rs1\[4\] i_rs1[4] _0994_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__mux2_1
X_6060_ reg_data\[6\]\[26\] _2207_ _2323_ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__and3_1
X_5011_ reg_data\[24\]\[9\] _1127_ _1130_ reg_data\[28\]\[9\] _1619_ vssd1 vssd1 vccd1
+ vccd1 _1620_ sky130_fd_sc_hd__a221o_1
X_6962_ _3336_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__clkbuf_1
X_9750_ clknet_leaf_16_i_clk _0894_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_9681_ clknet_leaf_21_i_clk _0825_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_5913_ reg_data\[18\]\[23\] _2422_ _2120_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__and3_1
X_6893_ reg_data\[2\]\[25\] _3181_ _3293_ vssd1 vssd1 vccd1 vccd1 _3299_ sky130_fd_sc_hd__mux2_1
X_8701_ _4277_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__clkbuf_1
X_5844_ reg_data\[3\]\[22\] _2421_ _2423_ _2424_ _2425_ vssd1 vssd1 vccd1 vccd1 _2426_
+ sky130_fd_sc_hd__a2111o_1
X_8632_ _3905_ reg_data\[12\]\[22\] _4238_ vssd1 vssd1 vccd1 vccd1 _4241_ sky130_fd_sc_hd__mux2_1
X_8563_ _4204_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__clkbuf_1
X_7514_ _3631_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__clkbuf_1
X_5775_ reg_data\[7\]\[21\] _1827_ _2356_ _2357_ _2358_ vssd1 vssd1 vccd1 vccd1 _2359_
+ sky130_fd_sc_hd__a2111o_1
X_8494_ _3903_ reg_data\[18\]\[21\] _4166_ vssd1 vssd1 vccd1 vccd1 _4168_ sky130_fd_sc_hd__mux2_1
X_4726_ _1163_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__clkbuf_4
X_7445_ _3256_ reg_data\[20\]\[26\] _3587_ vssd1 vssd1 vccd1 vccd1 _3594_ sky130_fd_sc_hd__mux2_1
X_4657_ reg_data\[25\]\[3\] _1141_ _1271_ _1274_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_
+ sky130_fd_sc_hd__a2111o_1
X_7376_ _3557_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__clkbuf_1
X_6327_ reg_data\[30\]\[31\] _2524_ _1056_ vssd1 vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__and3_1
X_4588_ reg_data\[23\]\[2\] _1206_ _1209_ reg_data\[19\]\[2\] vssd1 vssd1 vccd1 vccd1
+ _1210_ sky130_fd_sc_hd__a22o_1
X_9115_ clknet_leaf_3_i_clk _0259_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6258_ reg_data\[23\]\[29\] _2440_ _2441_ reg_data\[19\]\[29\] vssd1 vssd1 vccd1
+ vccd1 _2826_ sky130_fd_sc_hd__a22o_1
X_9046_ clknet_leaf_38_i_clk _0190_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6189_ reg_data\[21\]\[28\] _1162_ _1510_ vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__and3_1
X_5209_ reg_data\[22\]\[12\] _1679_ _1622_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__and3_1
X_9879_ clknet_leaf_49_i_clk _0949_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5560_ reg_data\[3\]\[18\] _1770_ _2148_ _2149_ _2150_ vssd1 vssd1 vccd1 vccd1 _2151_
+ sky130_fd_sc_hd__a2111o_1
X_5491_ reg_data\[22\]\[17\] _1536_ _1651_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__and3_1
X_4511_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__clkbuf_4
X_7230_ reg_data\[6\]\[21\] _3173_ _3478_ vssd1 vssd1 vccd1 vccd1 _3480_ sky130_fd_sc_hd__mux2_1
X_4442_ reg_data\[18\]\[2\] _1062_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__and3_1
X_4373_ i_rs2[0] i_rs2[1] i_rs_valid vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__o21a_1
X_7161_ _3443_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__clkbuf_1
X_6112_ reg_data\[30\]\[27\] _2204_ _1254_ vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__and3_1
X_7092_ _3406_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__clkbuf_1
X_6043_ reg_data\[2\]\[25\] _2443_ _2507_ _2508_ reg_data\[11\]\[25\] vssd1 vssd1
+ vccd1 vccd1 _2619_ sky130_fd_sc_hd__a32o_1
X_7994_ _3895_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__clkbuf_1
X_9802_ clknet_leaf_54_i_clk rdata1\[18\] vssd1 vssd1 vccd1 vccd1 r_data1\[18\] sky130_fd_sc_hd__dfxtp_1
X_6945_ _3327_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__clkbuf_1
X_9733_ clknet_leaf_65_i_clk _0877_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6876_ reg_data\[2\]\[17\] _3164_ _3282_ vssd1 vssd1 vccd1 vccd1 _3290_ sky130_fd_sc_hd__mux2_1
X_9664_ clknet_leaf_3_i_clk _0808_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_5827_ _1129_ vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__clkbuf_4
X_9595_ clknet_leaf_71_i_clk _0739_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_8615_ _3888_ reg_data\[12\]\[14\] _4227_ vssd1 vssd1 vccd1 vccd1 _4232_ sky130_fd_sc_hd__mux2_1
X_8546_ _4195_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__clkbuf_1
X_5758_ _2333_ _2338_ _2340_ _2342_ vssd1 vssd1 vccd1 vccd1 _2343_ sky130_fd_sc_hd__or4_1
X_4709_ reg_data\[2\]\[4\] _1103_ _1104_ _1106_ reg_data\[11\]\[4\] vssd1 vssd1 vccd1
+ vccd1 _1328_ sky130_fd_sc_hd__a32o_1
X_8477_ _3886_ reg_data\[18\]\[13\] _4155_ vssd1 vssd1 vccd1 vccd1 _4159_ sky130_fd_sc_hd__mux2_1
X_7428_ _3239_ reg_data\[20\]\[18\] _3576_ vssd1 vssd1 vccd1 vccd1 _3585_ sky130_fd_sc_hd__mux2_1
X_5689_ reg_data\[23\]\[20\] _1787_ _1788_ reg_data\[19\]\[20\] vssd1 vssd1 vccd1
+ vccd1 _2276_ sky130_fd_sc_hd__a22o_1
X_7359_ _3548_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__clkbuf_1
X_9029_ clknet_leaf_51_i_clk _0173_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6730_ reg_data\[4\]\[31\] _3193_ _3128_ vssd1 vssd1 vccd1 vccd1 _3194_ sky130_fd_sc_hd__mux2_1
X_4991_ _1071_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__clkbuf_4
X_6661_ i_data[9] vssd1 vssd1 vccd1 vccd1 _3147_ sky130_fd_sc_hd__buf_2
X_5612_ reg_data\[25\]\[19\] _1764_ _2198_ _2199_ _2200_ vssd1 vssd1 vccd1 vccd1 _2201_
+ sky130_fd_sc_hd__a2111o_1
X_9380_ clknet_leaf_59_i_clk _0524_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8400_ _3877_ reg_data\[17\]\[9\] _4108_ vssd1 vssd1 vccd1 vccd1 _4118_ sky130_fd_sc_hd__mux2_1
X_6592_ r_data2\[17\] _3094_ vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__and2_1
X_5543_ reg_data\[2\]\[17\] _1837_ _1901_ _1902_ reg_data\[11\]\[17\] vssd1 vssd1
+ vccd1 vccd1 _2135_ sky130_fd_sc_hd__a32o_1
X_8331_ _4081_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__clkbuf_1
X_8262_ _4044_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__clkbuf_1
X_5474_ reg_data\[5\]\[16\] _1824_ _1954_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__and3_1
X_4425_ _1047_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__clkbuf_4
X_7213_ reg_data\[6\]\[13\] _3156_ _3467_ vssd1 vssd1 vccd1 vccd1 _3471_ sky130_fd_sc_hd__mux2_1
X_8193_ _3875_ reg_data\[14\]\[8\] _3999_ vssd1 vssd1 vccd1 vccd1 _4008_ sky130_fd_sc_hd__mux2_1
X_7144_ _3434_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__clkbuf_1
X_7075_ _3397_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
X_6026_ reg_data\[21\]\[25\] _2489_ _1943_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__and3_1
X_7977_ i_data[12] vssd1 vssd1 vccd1 vccd1 _3884_ sky130_fd_sc_hd__buf_2
X_9716_ clknet_leaf_35_i_clk _0860_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6928_ _3318_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__clkbuf_1
X_9647_ clknet_leaf_30_i_clk _0791_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6859_ reg_data\[2\]\[9\] _3147_ _3271_ vssd1 vssd1 vccd1 vccd1 _3281_ sky130_fd_sc_hd__mux2_1
X_9578_ clknet_leaf_56_i_clk _0722_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8529_ _4186_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__clkbuf_1
X_5190_ _1108_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__clkbuf_4
X_7900_ _3837_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__clkbuf_1
X_8880_ clknet_leaf_23_i_clk _0024_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_7831_ _3800_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__clkbuf_1
X_4974_ reg_data\[1\]\[8\] _1298_ _1299_ reg_data\[15\]\[8\] vssd1 vssd1 vccd1 vccd1
+ _1584_ sky130_fd_sc_hd__a22o_1
X_7762_ _3229_ reg_data\[26\]\[13\] _3760_ vssd1 vssd1 vccd1 vccd1 _3764_ sky130_fd_sc_hd__mux2_1
X_6713_ _3182_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__clkbuf_1
X_7693_ _3727_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__clkbuf_1
X_9501_ clknet_leaf_4_i_clk _0645_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_9432_ clknet_leaf_69_i_clk _0576_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6644_ reg_data\[4\]\[3\] _3135_ _3129_ vssd1 vssd1 vccd1 vccd1 _3136_ sky130_fd_sc_hd__mux2_1
X_9363_ clknet_leaf_35_i_clk _0507_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6575_ r_data2\[9\] _3083_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__and2_1
X_9294_ clknet_leaf_39_i_clk _0438_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_5526_ reg_data\[17\]\[17\] _2117_ _1275_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__and3_1
X_8314_ _3857_ reg_data\[16\]\[0\] _4072_ vssd1 vssd1 vccd1 vccd1 _4073_ sky130_fd_sc_hd__mux2_1
X_8245_ _3857_ reg_data\[15\]\[0\] _4035_ vssd1 vssd1 vccd1 vccd1 _4036_ sky130_fd_sc_hd__mux2_1
X_5457_ reg_data\[8\]\[16\] _1797_ _1798_ reg_data\[10\]\[16\] _2051_ vssd1 vssd1
+ vccd1 vccd1 _2052_ sky130_fd_sc_hd__a221o_1
X_4408_ i_rs_valid rs1\[3\] vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__nor2_1
X_8176_ _3998_ vssd1 vssd1 vccd1 vccd1 _3999_ sky130_fd_sc_hd__clkbuf_4
X_5388_ reg_data\[13\]\[15\] _1867_ _1087_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__and3_1
X_7127_ _3425_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
X_7058_ _3388_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__clkbuf_1
X_6009_ reg_data\[0\]\[25\] _2381_ _2583_ _2584_ _2585_ vssd1 vssd1 vccd1 vccd1 _2586_
+ sky130_fd_sc_hd__a2111o_1
X_4690_ reg_data\[17\]\[4\] _1046_ _1108_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__and3_1
X_6360_ reg_data\[5\]\[31\] _2430_ _1338_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__and3_1
X_5311_ reg_data\[24\]\[13\] _1847_ _1848_ reg_data\[28\]\[13\] _1910_ vssd1 vssd1
+ vccd1 vccd1 _1911_ sky130_fd_sc_hd__a221o_1
X_8030_ _3919_ reg_data\[9\]\[29\] _3901_ vssd1 vssd1 vccd1 vccd1 _3920_ sky130_fd_sc_hd__mux2_1
X_6291_ reg_data\[26\]\[30\] _2411_ _2412_ reg_data\[29\]\[30\] vssd1 vssd1 vccd1
+ vccd1 _2858_ sky130_fd_sc_hd__a22o_1
X_5242_ _1220_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__clkbuf_4
X_5173_ reg_data\[6\]\[12\] _1600_ _1716_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__and3_1
X_8932_ clknet_leaf_60_i_clk _0076_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8863_ clknet_leaf_2_i_clk _0007_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_7814_ _3791_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__clkbuf_1
X_8794_ reg_data\[11\]\[2\] i_data[2] _4324_ vssd1 vssd1 vccd1 vccd1 _4327_ sky130_fd_sc_hd__mux2_1
X_7745_ _3212_ reg_data\[26\]\[5\] _3749_ vssd1 vssd1 vccd1 vccd1 _3755_ sky130_fd_sc_hd__mux2_1
X_4957_ reg_data\[18\]\[8\] _1159_ _1513_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__and3_1
X_4888_ reg_data\[27\]\[7\] _1096_ _1498_ _1499_ _1500_ vssd1 vssd1 vccd1 vccd1 _1501_
+ sky130_fd_sc_hd__a2111o_1
X_7676_ _3718_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__clkbuf_1
X_9415_ clknet_leaf_53_i_clk _0559_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6627_ i_rd[3] _3119_ vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__or2_1
X_9346_ clknet_leaf_59_i_clk _0490_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6558_ _3084_ vssd1 vssd1 vccd1 vccd1 o_data2[0] sky130_fd_sc_hd__buf_2
X_5509_ _1086_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__clkbuf_4
X_9277_ clknet_leaf_69_i_clk _0421_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6489_ _3047_ vssd1 vssd1 vccd1 vccd1 o_data1[0] sky130_fd_sc_hd__buf_2
X_8228_ _4026_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__clkbuf_1
X_8159_ _3909_ reg_data\[13\]\[24\] _3985_ vssd1 vssd1 vccd1 vccd1 _3990_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_7_i_clk clknet_3_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5860_ reg_data\[23\]\[22\] _2440_ _2441_ reg_data\[19\]\[22\] vssd1 vssd1 vccd1
+ vccd1 _2442_ sky130_fd_sc_hd__a22o_1
X_4811_ reg_data\[17\]\[6\] _1042_ _1238_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__and3_1
X_5791_ reg_data\[21\]\[22\] _2086_ _2087_ vssd1 vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__and3_1
X_4742_ reg_data\[1\]\[4\] _1298_ _1299_ reg_data\[15\]\[4\] vssd1 vssd1 vccd1 vccd1
+ _1360_ sky130_fd_sc_hd__a22o_1
X_7530_ reg_data\[23\]\[0\] _3118_ _3640_ vssd1 vssd1 vccd1 vccd1 _3641_ sky130_fd_sc_hd__mux2_1
X_7461_ _3195_ reg_data\[21\]\[0\] _3603_ vssd1 vssd1 vccd1 vccd1 _3604_ sky130_fd_sc_hd__mux2_1
X_4673_ _1277_ _1281_ _1287_ _1292_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__or4_1
X_9200_ clknet_leaf_22_i_clk _0344_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6412_ reg_data\[6\]\[0\] _2555_ _1270_ vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__and3_1
X_7392_ _3566_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__clkbuf_1
X_6343_ reg_data\[16\]\[31\] _2405_ _2406_ reg_data\[9\]\[31\] vssd1 vssd1 vccd1 vccd1
+ _2908_ sky130_fd_sc_hd__a22o_1
X_9131_ clknet_leaf_27_i_clk _0275_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6274_ reg_data\[20\]\[30\] _1046_ _2035_ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__and3_1
X_9062_ clknet_leaf_45_i_clk _0206_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8013_ _3908_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__clkbuf_1
X_5225_ _1184_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__clkbuf_4
X_5156_ reg_data\[8\]\[11\] _1214_ _1217_ reg_data\[10\]\[11\] _1759_ vssd1 vssd1
+ vccd1 vccd1 _1760_ sky130_fd_sc_hd__a221o_1
X_5087_ _1171_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__buf_2
X_8915_ clknet_leaf_21_i_clk _0059_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_9895_ clknet_leaf_77_i_clk _0965_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_8846_ reg_data\[11\]\[27\] i_data[27] _4346_ vssd1 vssd1 vccd1 vccd1 _4354_ sky130_fd_sc_hd__mux2_1
X_8777_ _4317_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__clkbuf_1
X_5989_ reg_data\[2\]\[24\] _2443_ _2507_ _2508_ reg_data\[11\]\[24\] vssd1 vssd1
+ vccd1 vccd1 _2567_ sky130_fd_sc_hd__a32o_1
X_7728_ _3745_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__clkbuf_1
X_7659_ _3262_ reg_data\[24\]\[29\] _3699_ vssd1 vssd1 vccd1 vccd1 _3709_ sky130_fd_sc_hd__mux2_1
X_9329_ clknet_leaf_22_i_clk _0473_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_5010_ reg_data\[26\]\[9\] _1132_ _1134_ reg_data\[29\]\[9\] vssd1 vssd1 vccd1 vccd1
+ _1619_ sky130_fd_sc_hd__a22o_1
X_6961_ _3252_ reg_data\[10\]\[24\] _3331_ vssd1 vssd1 vccd1 vccd1 _3336_ sky130_fd_sc_hd__mux2_1
X_8700_ reg_data\[19\]\[22\] _3175_ _4274_ vssd1 vssd1 vccd1 vccd1 _4277_ sky130_fd_sc_hd__mux2_1
X_9680_ clknet_leaf_18_i_clk _0824_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_5912_ reg_data\[25\]\[23\] _2416_ _2488_ _2490_ _2491_ vssd1 vssd1 vccd1 vccd1 _2492_
+ sky130_fd_sc_hd__a2111o_1
X_6892_ _3298_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__clkbuf_1
X_5843_ reg_data\[20\]\[22\] _2234_ _1743_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__and3_1
X_8631_ _4240_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__clkbuf_1
X_8562_ reg_data\[1\]\[21\] _3173_ _4202_ vssd1 vssd1 vccd1 vccd1 _4204_ sky130_fd_sc_hd__mux2_1
X_7513_ _3254_ reg_data\[21\]\[25\] _3625_ vssd1 vssd1 vccd1 vccd1 _3631_ sky130_fd_sc_hd__mux2_1
X_5774_ reg_data\[12\]\[21\] _1960_ _2016_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__and3_1
X_8493_ _4167_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__clkbuf_1
X_4725_ reg_data\[20\]\[4\] _1162_ _1342_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__and3_1
X_7444_ _3593_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__clkbuf_1
X_4656_ reg_data\[17\]\[3\] _1150_ _1275_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__and3_1
X_7375_ reg_data\[3\]\[25\] _3181_ _3551_ vssd1 vssd1 vccd1 vccd1 _3557_ sky130_fd_sc_hd__mux2_1
X_4587_ _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__buf_4
X_6326_ reg_data\[18\]\[31\] _1039_ _1063_ vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__and3_1
X_9114_ clknet_leaf_12_i_clk _0258_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6257_ _2812_ _2816_ _2820_ _2824_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__or4_4
X_9045_ clknet_leaf_37_i_clk _0189_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6188_ reg_data\[17\]\[28\] _2489_ _1395_ vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__and3_1
X_5208_ _1140_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_72_i_clk clknet_3_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5139_ _1160_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__clkbuf_4
X_9878_ clknet_leaf_49_i_clk _0948_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8829_ reg_data\[11\]\[19\] i_data[19] _4335_ vssd1 vssd1 vccd1 vccd1 _4345_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_i_clk clknet_3_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_25_i_clk clknet_3_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4510_ _1058_ _1086_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__and2_4
X_5490_ _2083_ vssd1 vssd1 vccd1 vccd1 rdata2\[16\] sky130_fd_sc_hd__clkbuf_1
X_4441_ _1063_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__buf_4
X_7160_ reg_data\[7\]\[20\] _3170_ _3442_ vssd1 vssd1 vccd1 vccd1 _3443_ sky130_fd_sc_hd__mux2_1
X_6111_ reg_data\[20\]\[27\] _2524_ _1059_ vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__and3_1
X_4372_ i_rs2[0] i_rs2[1] vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__nand2_1
X_7091_ _3243_ reg_data\[8\]\[20\] _3405_ vssd1 vssd1 vccd1 vccd1 _3406_ sky130_fd_sc_hd__mux2_1
X_6042_ reg_data\[23\]\[25\] _2440_ _2441_ reg_data\[19\]\[25\] vssd1 vssd1 vccd1
+ vccd1 _2618_ sky130_fd_sc_hd__a22o_1
X_9801_ clknet_leaf_54_i_clk rdata1\[17\] vssd1 vssd1 vccd1 vccd1 r_data1\[17\] sky130_fd_sc_hd__dfxtp_1
X_7993_ _3894_ reg_data\[9\]\[17\] _3880_ vssd1 vssd1 vccd1 vccd1 _3895_ sky130_fd_sc_hd__mux2_1
X_6944_ _3235_ reg_data\[10\]\[16\] _3320_ vssd1 vssd1 vccd1 vccd1 _3327_ sky130_fd_sc_hd__mux2_1
X_9732_ clknet_leaf_65_i_clk _0876_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_9663_ clknet_leaf_5_i_clk _0807_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6875_ _3289_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__clkbuf_1
X_8614_ _4231_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__clkbuf_1
X_5826_ _1126_ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__clkbuf_4
X_9594_ clknet_leaf_70_i_clk _0738_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8545_ reg_data\[1\]\[13\] _3156_ _4191_ vssd1 vssd1 vccd1 vccd1 _4195_ sky130_fd_sc_hd__mux2_1
X_5757_ reg_data\[24\]\[21\] _1803_ _1804_ reg_data\[28\]\[21\] _2341_ vssd1 vssd1
+ vccd1 vccd1 _2342_ sky130_fd_sc_hd__a221o_1
X_4708_ reg_data\[23\]\[4\] _1099_ _1101_ reg_data\[19\]\[4\] vssd1 vssd1 vccd1 vccd1
+ _1327_ sky130_fd_sc_hd__a22o_1
X_8476_ _4158_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__clkbuf_1
X_5688_ _2260_ _2265_ _2269_ _2274_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__or4_2
X_7427_ _3584_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__clkbuf_1
X_4639_ _1242_ _1246_ _1252_ _1259_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__or4_1
X_7358_ reg_data\[3\]\[17\] _3164_ _3540_ vssd1 vssd1 vccd1 vccd1 _3548_ sky130_fd_sc_hd__mux2_1
X_6309_ reg_data\[12\]\[30\] _2562_ _1289_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__and3_1
X_7289_ _3511_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__clkbuf_1
X_9028_ clknet_leaf_62_i_clk _0172_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_4990_ reg_data\[3\]\[9\] _1054_ _1595_ _1596_ _1598_ vssd1 vssd1 vccd1 vccd1 _1599_
+ sky130_fd_sc_hd__a2111o_1
X_6660_ _3146_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__clkbuf_1
X_5611_ reg_data\[17\]\[19\] _2086_ _1238_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__and3_1
X_6591_ _3101_ vssd1 vssd1 vccd1 vccd1 o_data2[16] sky130_fd_sc_hd__buf_2
X_8330_ _3875_ reg_data\[16\]\[8\] _4072_ vssd1 vssd1 vccd1 vccd1 _4081_ sky130_fd_sc_hd__mux2_1
X_5542_ reg_data\[23\]\[17\] _1834_ _1835_ reg_data\[19\]\[17\] vssd1 vssd1 vccd1
+ vccd1 _2134_ sky130_fd_sc_hd__a22o_1
X_8261_ _3875_ reg_data\[15\]\[8\] _4035_ vssd1 vssd1 vccd1 vccd1 _4044_ sky130_fd_sc_hd__mux2_1
X_5473_ reg_data\[4\]\[16\] _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__and3_1
X_4424_ _1025_ _1033_ rs1_mux\[2\] _1015_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__and4b_4
X_7212_ _3470_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_1
X_8192_ _4007_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__clkbuf_1
X_7143_ reg_data\[7\]\[12\] _3154_ _3431_ vssd1 vssd1 vccd1 vccd1 _3434_ sky130_fd_sc_hd__mux2_1
X_7074_ _3227_ reg_data\[8\]\[12\] _3394_ vssd1 vssd1 vccd1 vccd1 _3397_ sky130_fd_sc_hd__mux2_1
X_6025_ reg_data\[22\]\[25\] _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__and3_1
X_9715_ clknet_leaf_35_i_clk _0859_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_7976_ _3883_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__clkbuf_1
X_6927_ _3218_ reg_data\[10\]\[8\] _3309_ vssd1 vssd1 vccd1 vccd1 _3318_ sky130_fd_sc_hd__mux2_1
X_9646_ clknet_leaf_29_i_clk _0790_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6858_ _3280_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__clkbuf_1
X_5809_ _1095_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__clkbuf_4
X_9577_ clknet_leaf_59_i_clk _0721_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_8528_ reg_data\[1\]\[5\] _3139_ _4180_ vssd1 vssd1 vccd1 vccd1 _4186_ sky130_fd_sc_hd__mux2_1
X_6789_ _3235_ reg_data\[22\]\[16\] _3223_ vssd1 vssd1 vccd1 vccd1 _3236_ sky130_fd_sc_hd__mux2_1
X_8459_ _4149_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__clkbuf_1
X_7830_ _3229_ reg_data\[27\]\[13\] _3796_ vssd1 vssd1 vccd1 vccd1 _3800_ sky130_fd_sc_hd__mux2_1
X_4973_ reg_data\[2\]\[8\] _1002_ _1295_ _1296_ reg_data\[11\]\[8\] vssd1 vssd1 vccd1
+ vccd1 _1583_ sky130_fd_sc_hd__a32o_1
X_7761_ _3763_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__clkbuf_1
X_6712_ reg_data\[4\]\[25\] _3181_ _3171_ vssd1 vssd1 vccd1 vccd1 _3182_ sky130_fd_sc_hd__mux2_1
X_7692_ _3227_ reg_data\[25\]\[12\] _3724_ vssd1 vssd1 vccd1 vccd1 _3727_ sky130_fd_sc_hd__mux2_1
X_9500_ clknet_leaf_11_i_clk _0644_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_9431_ clknet_leaf_43_i_clk _0575_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6643_ i_data[3] vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__buf_2
X_9362_ clknet_leaf_34_i_clk _0506_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6574_ _3092_ vssd1 vssd1 vccd1 vccd1 o_data2[8] sky130_fd_sc_hd__buf_2
X_5525_ _1138_ vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__buf_4
X_8313_ _4071_ vssd1 vssd1 vccd1 vccd1 _4072_ sky130_fd_sc_hd__buf_4
X_9293_ clknet_leaf_49_i_clk _0437_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_8244_ _4034_ vssd1 vssd1 vccd1 vccd1 _4035_ sky130_fd_sc_hd__buf_4
X_5456_ reg_data\[16\]\[16\] _1799_ _1800_ reg_data\[9\]\[16\] vssd1 vssd1 vccd1 vccd1
+ _2051_ sky130_fd_sc_hd__a22o_1
X_4407_ i_rs1[0] i_rs1[2] i_rs1[1] i_rs1[3] vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__o31ai_1
X_8175_ _3200_ _3961_ vssd1 vssd1 vccd1 vccd1 _3998_ sky130_fd_sc_hd__nand2_4
X_5387_ reg_data\[0\]\[15\] _1775_ _1981_ _1982_ _1983_ vssd1 vssd1 vccd1 vccd1 _1984_
+ sky130_fd_sc_hd__a2111o_1
X_7126_ reg_data\[7\]\[4\] _3137_ _3420_ vssd1 vssd1 vccd1 vccd1 _3425_ sky130_fd_sc_hd__mux2_1
X_7057_ _3210_ reg_data\[8\]\[4\] _3383_ vssd1 vssd1 vccd1 vccd1 _3388_ sky130_fd_sc_hd__mux2_1
X_6008_ reg_data\[5\]\[25\] _2097_ _2530_ vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__and3_1
X_7959_ _3871_ reg_data\[9\]\[6\] _3859_ vssd1 vssd1 vccd1 vccd1 _3872_ sky130_fd_sc_hd__mux2_1
X_9629_ clknet_leaf_7_i_clk _0773_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6290_ reg_data\[8\]\[30\] _2403_ _2404_ reg_data\[10\]\[30\] _2856_ vssd1 vssd1
+ vccd1 vccd1 _2857_ sky130_fd_sc_hd__a221o_1
X_5310_ reg_data\[26\]\[13\] _1849_ _1850_ reg_data\[29\]\[13\] vssd1 vssd1 vccd1
+ vccd1 _1910_ sky130_fd_sc_hd__a22o_1
X_5241_ _1218_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__clkbuf_4
X_5172_ _1069_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__buf_4
X_8931_ clknet_leaf_61_i_clk _0075_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8862_ clknet_leaf_3_i_clk _0006_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_7813_ _3212_ reg_data\[27\]\[5\] _3785_ vssd1 vssd1 vccd1 vccd1 _3791_ sky130_fd_sc_hd__mux2_1
X_8793_ _4326_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__clkbuf_1
X_7744_ _3754_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__clkbuf_1
X_4956_ reg_data\[25\]\[8\] _1141_ _1563_ _1564_ _1565_ vssd1 vssd1 vccd1 vccd1 _1566_
+ sky130_fd_sc_hd__a2111o_1
X_4887_ reg_data\[1\]\[7\] _1022_ _1109_ _1111_ reg_data\[15\]\[7\] vssd1 vssd1 vccd1
+ vccd1 _1500_ sky130_fd_sc_hd__a32o_1
X_7675_ _3210_ reg_data\[25\]\[4\] _3713_ vssd1 vssd1 vccd1 vccd1 _3718_ sky130_fd_sc_hd__mux2_1
X_6626_ _3119_ _3120_ vssd1 vssd1 vccd1 vccd1 _3121_ sky130_fd_sc_hd__and2_1
X_9414_ clknet_leaf_54_i_clk _0558_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_9345_ clknet_leaf_72_i_clk _0489_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6557_ r_data2\[0\] _3083_ vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__and2_1
X_5508_ reg_data\[12\]\[17\] _1986_ _1606_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__and3_1
X_9276_ clknet_leaf_71_i_clk _0420_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6488_ r_data1\[0\] _3046_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__and2_1
X_8227_ _3909_ reg_data\[14\]\[24\] _4021_ vssd1 vssd1 vccd1 vccd1 _4026_ sky130_fd_sc_hd__mux2_1
X_5439_ reg_data\[30\]\[16\] _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__and3_1
X_8158_ _3989_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__clkbuf_1
X_7109_ _3262_ reg_data\[8\]\[29\] _3405_ vssd1 vssd1 vccd1 vccd1 _3415_ sky130_fd_sc_hd__mux2_1
X_8089_ _3952_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__clkbuf_1
X_4810_ reg_data\[22\]\[6\] _1039_ _1236_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__and3_1
X_5790_ reg_data\[17\]\[22\] _2372_ _1708_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__and3_1
X_4741_ reg_data\[2\]\[4\] _1002_ _1295_ _1296_ reg_data\[11\]\[4\] vssd1 vssd1 vccd1
+ vccd1 _1359_ sky130_fd_sc_hd__a32o_1
X_7460_ _3602_ vssd1 vssd1 vccd1 vccd1 _3603_ sky130_fd_sc_hd__buf_4
X_4672_ reg_data\[7\]\[3\] _1185_ _1288_ _1290_ _1291_ vssd1 vssd1 vccd1 vccd1 _1292_
+ sky130_fd_sc_hd__a2111o_1
X_6411_ reg_data\[3\]\[0\] _1157_ _2970_ _2971_ _2972_ vssd1 vssd1 vccd1 vccd1 _2973_
+ sky130_fd_sc_hd__a2111o_1
X_9130_ clknet_leaf_43_i_clk _0274_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_7391_ _3195_ reg_data\[20\]\[0\] _3565_ vssd1 vssd1 vccd1 vccd1 _3566_ sky130_fd_sc_hd__mux2_1
X_6342_ reg_data\[27\]\[31\] _2392_ _2904_ _2905_ _2906_ vssd1 vssd1 vccd1 vccd1 _2907_
+ sky130_fd_sc_hd__a2111o_1
X_6273_ reg_data\[30\]\[30\] _2524_ _1919_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__and3_1
X_9061_ clknet_leaf_63_i_clk _0205_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8012_ _3907_ reg_data\[9\]\[23\] _3901_ vssd1 vssd1 vccd1 vccd1 _3908_ sky130_fd_sc_hd__mux2_1
X_5224_ reg_data\[0\]\[12\] _1821_ _1822_ _1823_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_
+ sky130_fd_sc_hd__a2111o_1
X_5155_ reg_data\[16\]\[11\] _1219_ _1221_ reg_data\[9\]\[11\] vssd1 vssd1 vccd1 vccd1
+ _1759_ sky130_fd_sc_hd__a22o_1
X_5086_ reg_data\[13\]\[10\] _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__and3_1
X_8914_ clknet_leaf_30_i_clk _0058_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_9894_ clknet_leaf_75_i_clk _0964_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_8845_ _4353_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__clkbuf_1
X_8776_ _3913_ reg_data\[29\]\[26\] _4310_ vssd1 vssd1 vccd1 vccd1 _4317_ sky130_fd_sc_hd__mux2_1
X_5988_ reg_data\[23\]\[24\] _2440_ _2441_ reg_data\[19\]\[24\] vssd1 vssd1 vccd1
+ vccd1 _2566_ sky130_fd_sc_hd__a22o_1
X_7727_ _3262_ reg_data\[25\]\[29\] _3735_ vssd1 vssd1 vccd1 vccd1 _3745_ sky130_fd_sc_hd__mux2_1
X_4939_ reg_data\[12\]\[8\] _1381_ _1128_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__and3_1
X_7658_ _3708_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__clkbuf_1
X_6609_ r_data2\[25\] _3105_ vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__and2_1
X_7589_ _3671_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__clkbuf_1
X_9328_ clknet_leaf_22_i_clk _0472_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_9259_ clknet_leaf_59_i_clk _0403_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6960_ _3335_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__clkbuf_1
X_5911_ reg_data\[21\]\[23\] _2117_ _1510_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__and3_1
X_6891_ reg_data\[2\]\[24\] _3179_ _3293_ vssd1 vssd1 vccd1 vccd1 _3298_ sky130_fd_sc_hd__mux2_1
X_5842_ reg_data\[30\]\[22\] _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__and3_1
X_8630_ _3903_ reg_data\[12\]\[21\] _4238_ vssd1 vssd1 vccd1 vccd1 _4240_ sky130_fd_sc_hd__mux2_1
X_5773_ reg_data\[14\]\[21\] _2301_ _1958_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__and3_1
X_8561_ _4203_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__clkbuf_1
X_7512_ _3630_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__clkbuf_1
X_4724_ _1160_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__clkbuf_4
X_8492_ _3900_ reg_data\[18\]\[20\] _4166_ vssd1 vssd1 vccd1 vccd1 _4167_ sky130_fd_sc_hd__mux2_1
X_7443_ _3254_ reg_data\[20\]\[25\] _3587_ vssd1 vssd1 vccd1 vccd1 _3593_ sky130_fd_sc_hd__mux2_1
X_4655_ _1147_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__clkbuf_4
X_7374_ _3556_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__clkbuf_1
X_4586_ _1207_ _1155_ _1156_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_6_i_clk clknet_3_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_6325_ reg_data\[25\]\[31\] _2370_ _2887_ _2888_ _2889_ vssd1 vssd1 vccd1 vccd1 _2890_
+ sky130_fd_sc_hd__a2111o_1
X_9113_ clknet_leaf_13_i_clk _0257_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_9044_ clknet_leaf_32_i_clk _0188_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6256_ reg_data\[7\]\[29\] _2433_ _2821_ _2822_ _2823_ vssd1 vssd1 vccd1 vccd1 _2824_
+ sky130_fd_sc_hd__a2111o_1
X_6187_ reg_data\[22\]\[28\] _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__and3_1
X_5207_ _1809_ vssd1 vssd1 vccd1 vccd1 rdata1\[12\] sky130_fd_sc_hd__clkbuf_1
X_5138_ reg_data\[30\]\[11\] _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__and3_1
X_5069_ reg_data\[26\]\[10\] _1132_ _1134_ reg_data\[29\]\[10\] vssd1 vssd1 vccd1
+ vccd1 _1676_ sky130_fd_sc_hd__a22o_1
X_9877_ clknet_leaf_59_i_clk _0947_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_8828_ _4344_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__clkbuf_1
X_8759_ _3896_ reg_data\[29\]\[18\] _4299_ vssd1 vssd1 vccd1 vccd1 _4308_ sky130_fd_sc_hd__mux2_1
X_4440_ rs1_mux\[0\] _1025_ _1030_ _1033_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__and4bb_2
X_6110_ reg_data\[18\]\[27\] _2261_ _1063_ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__and3_1
X_4371_ _1002_ vssd1 vssd1 vccd1 vccd1 rs2_mux\[4\] sky130_fd_sc_hd__inv_2
X_7090_ _3382_ vssd1 vssd1 vccd1 vccd1 _3405_ sky130_fd_sc_hd__buf_4
X_6041_ _2604_ _2608_ _2612_ _2616_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__or4_2
X_9800_ clknet_leaf_54_i_clk rdata1\[16\] vssd1 vssd1 vccd1 vccd1 r_data1\[16\] sky130_fd_sc_hd__dfxtp_1
X_7992_ i_data[17] vssd1 vssd1 vccd1 vccd1 _3894_ sky130_fd_sc_hd__clkbuf_4
X_6943_ _3326_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__clkbuf_1
X_9731_ clknet_leaf_7_i_clk _0875_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6874_ reg_data\[2\]\[16\] _3162_ _3282_ vssd1 vssd1 vccd1 vccd1 _3289_ sky130_fd_sc_hd__mux2_1
X_9662_ clknet_leaf_3_i_clk _0806_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_5825_ reg_data\[8\]\[22\] _2403_ _2404_ reg_data\[10\]\[22\] _2407_ vssd1 vssd1
+ vccd1 vccd1 _2408_ sky130_fd_sc_hd__a221o_1
X_8613_ _3886_ reg_data\[12\]\[13\] _4227_ vssd1 vssd1 vccd1 vccd1 _4231_ sky130_fd_sc_hd__mux2_1
X_9593_ clknet_leaf_67_i_clk _0737_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8544_ _4194_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__clkbuf_1
X_5756_ reg_data\[26\]\[21\] _1805_ _1806_ reg_data\[29\]\[21\] vssd1 vssd1 vccd1
+ vccd1 _2341_ sky130_fd_sc_hd__a22o_1
X_5687_ reg_data\[7\]\[20\] _1780_ _2270_ _2272_ _2273_ vssd1 vssd1 vccd1 vccd1 _2274_
+ sky130_fd_sc_hd__a2111o_1
X_8475_ _3884_ reg_data\[18\]\[12\] _4155_ vssd1 vssd1 vccd1 vccd1 _4158_ sky130_fd_sc_hd__mux2_1
X_4707_ _1310_ _1317_ _1321_ _1325_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__or4_1
X_4638_ reg_data\[7\]\[3\] _1081_ _1255_ _1256_ _1258_ vssd1 vssd1 vccd1 vccd1 _1259_
+ sky130_fd_sc_hd__a2111o_1
X_7426_ _3237_ reg_data\[20\]\[17\] _3576_ vssd1 vssd1 vccd1 vccd1 _3584_ sky130_fd_sc_hd__mux2_1
X_4569_ _1190_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__clkbuf_4
X_7357_ _3547_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__clkbuf_1
X_6308_ reg_data\[14\]\[30\] _1186_ _1344_ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__and3_1
X_7288_ reg_data\[5\]\[16\] _3162_ _3504_ vssd1 vssd1 vccd1 vccd1 _3511_ sky130_fd_sc_hd__mux2_1
X_6239_ _2799_ _2803_ _2805_ _2807_ vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__or4_1
X_9027_ clknet_leaf_59_i_clk _0171_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_5610_ reg_data\[21\]\[19\] _1766_ _1043_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_71_i_clk clknet_3_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_6590_ r_data2\[16\] _3094_ vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__and2_1
X_5541_ _2119_ _2124_ _2128_ _2132_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__or4_1
X_8260_ _4043_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__clkbuf_1
X_5472_ _1160_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__buf_2
X_7211_ reg_data\[6\]\[12\] _3154_ _3467_ vssd1 vssd1 vccd1 vccd1 _3470_ sky130_fd_sc_hd__mux2_1
X_4423_ _1034_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__buf_2
X_8191_ _3873_ reg_data\[14\]\[7\] _3999_ vssd1 vssd1 vccd1 vccd1 _4007_ sky130_fd_sc_hd__mux2_1
X_7142_ _3433_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__clkbuf_1
X_7073_ _3396_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
X_6024_ _2600_ vssd1 vssd1 vccd1 vccd1 rdata1\[25\] sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_24_i_clk clknet_3_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_7975_ _3882_ reg_data\[9\]\[11\] _3880_ vssd1 vssd1 vccd1 vccd1 _3883_ sky130_fd_sc_hd__mux2_1
X_9714_ clknet_leaf_35_i_clk _0858_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6926_ _3317_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__clkbuf_1
X_9645_ clknet_leaf_43_i_clk _0789_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6857_ reg_data\[2\]\[8\] _3145_ _3271_ vssd1 vssd1 vccd1 vccd1 _3280_ sky130_fd_sc_hd__mux2_1
X_5808_ _2375_ _2380_ _2385_ _2390_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_39_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_9576_ clknet_leaf_56_i_clk _0720_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6788_ i_data[16] vssd1 vssd1 vccd1 vccd1 _3235_ sky130_fd_sc_hd__buf_2
X_5739_ reg_data\[6\]\[21\] _2207_ _2323_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__and3_1
X_8527_ _4185_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__clkbuf_1
X_8458_ _3867_ reg_data\[18\]\[4\] _4144_ vssd1 vssd1 vccd1 vccd1 _4149_ sky130_fd_sc_hd__mux2_1
X_7409_ _3220_ reg_data\[20\]\[9\] _3565_ vssd1 vssd1 vccd1 vccd1 _3575_ sky130_fd_sc_hd__mux2_1
X_8389_ _4112_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__clkbuf_1
X_4972_ reg_data\[23\]\[8\] _1206_ _1209_ reg_data\[19\]\[8\] vssd1 vssd1 vccd1 vccd1
+ _1582_ sky130_fd_sc_hd__a22o_1
X_7760_ _3227_ reg_data\[26\]\[12\] _3760_ vssd1 vssd1 vccd1 vccd1 _3763_ sky130_fd_sc_hd__mux2_1
X_6711_ i_data[25] vssd1 vssd1 vccd1 vccd1 _3181_ sky130_fd_sc_hd__buf_4
X_7691_ _3726_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__clkbuf_1
X_9430_ clknet_leaf_38_i_clk _0574_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6642_ _3134_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__clkbuf_1
X_9361_ clknet_leaf_35_i_clk _0505_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_8312_ _3381_ _4070_ vssd1 vssd1 vccd1 vccd1 _4071_ sky130_fd_sc_hd__nand2_4
X_6573_ r_data2\[8\] _3083_ vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__and2_1
X_5524_ reg_data\[21\]\[17\] _1883_ _1943_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__and3_1
X_9292_ clknet_leaf_50_i_clk _0436_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8243_ _3638_ _3961_ vssd1 vssd1 vccd1 vccd1 _4034_ sky130_fd_sc_hd__nand2_4
X_5455_ reg_data\[27\]\[16\] _1786_ _2047_ _2048_ _2049_ vssd1 vssd1 vccd1 vccd1 _2050_
+ sky130_fd_sc_hd__a2111o_1
X_4406_ _1030_ vssd1 vssd1 vccd1 vccd1 rs1_mux\[2\] sky130_fd_sc_hd__clkinv_2
X_8174_ _3997_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__clkbuf_1
X_7125_ _3424_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
X_5386_ reg_data\[5\]\[15\] _1490_ _1925_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__and3_1
X_7056_ _3387_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__clkbuf_1
X_6007_ reg_data\[4\]\[25\] _2325_ _2469_ vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__and3_1
X_7958_ i_data[6] vssd1 vssd1 vccd1 vccd1 _3871_ sky130_fd_sc_hd__clkbuf_4
X_6909_ _3200_ _3307_ vssd1 vssd1 vccd1 vccd1 _3308_ sky130_fd_sc_hd__nand2_4
X_7889_ _3831_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__clkbuf_1
X_9628_ clknet_leaf_7_i_clk _0772_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_9559_ clknet_leaf_13_i_clk _0703_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5240_ _1216_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__buf_2
X_5171_ reg_data\[3\]\[12\] _1770_ _1771_ _1772_ _1773_ vssd1 vssd1 vccd1 vccd1 _1774_
+ sky130_fd_sc_hd__a2111o_1
X_8930_ clknet_leaf_60_i_clk _0074_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8861_ clknet_leaf_3_i_clk _0005_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_7812_ _3790_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__clkbuf_1
X_8792_ reg_data\[11\]\[1\] i_data[1] _4324_ vssd1 vssd1 vccd1 vccd1 _4326_ sky130_fd_sc_hd__mux2_1
X_7743_ _3210_ reg_data\[26\]\[4\] _3749_ vssd1 vssd1 vccd1 vccd1 _3754_ sky130_fd_sc_hd__mux2_1
X_4955_ reg_data\[21\]\[8\] _1509_ _1510_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__and3_1
X_4886_ reg_data\[2\]\[7\] _1103_ _1104_ _1106_ reg_data\[11\]\[7\] vssd1 vssd1 vccd1
+ vccd1 _1499_ sky130_fd_sc_hd__a32o_1
X_7674_ _3717_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__clkbuf_1
X_9413_ clknet_leaf_52_i_clk _0557_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6625_ i_rd[0] i_rd[1] i_rd[2] vssd1 vssd1 vccd1 vccd1 _3120_ sky130_fd_sc_hd__o21ai_1
X_9344_ clknet_leaf_70_i_clk _0488_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6556_ _3082_ vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__dlymetal6s2s_1
X_5507_ reg_data\[14\]\[17\] _1867_ _1379_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__and3_1
X_9275_ clknet_leaf_70_i_clk _0419_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_8226_ _4025_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__clkbuf_1
X_6487_ _3045_ vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__clkbuf_2
X_5438_ reg_data\[18\]\[16\] _1656_ _1483_ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__and3_1
X_8157_ _3907_ reg_data\[13\]\[23\] _3985_ vssd1 vssd1 vccd1 vccd1 _3989_ sky130_fd_sc_hd__mux2_1
X_5369_ reg_data\[27\]\[14\] _1833_ _1964_ _1965_ _1966_ vssd1 vssd1 vccd1 vccd1 _1967_
+ sky130_fd_sc_hd__a2111o_1
X_8088_ _3907_ reg_data\[30\]\[23\] _3948_ vssd1 vssd1 vccd1 vccd1 _3952_ sky130_fd_sc_hd__mux2_1
X_7108_ _3414_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
X_7039_ reg_data\[0\]\[29\] _3189_ _3367_ vssd1 vssd1 vccd1 vccd1 _3377_ sky130_fd_sc_hd__mux2_1
X_4740_ reg_data\[23\]\[4\] _1206_ _1209_ reg_data\[19\]\[4\] vssd1 vssd1 vccd1 vccd1
+ _1358_ sky130_fd_sc_hd__a22o_1
X_4671_ reg_data\[13\]\[3\] _1001_ _1191_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__and3_1
X_6410_ reg_data\[20\]\[0\] _1150_ _1283_ vssd1 vssd1 vccd1 vccd1 _2972_ sky130_fd_sc_hd__and3_1
X_7390_ _3564_ vssd1 vssd1 vccd1 vccd1 _3565_ sky130_fd_sc_hd__buf_4
X_6341_ reg_data\[1\]\[31\] _1103_ _2399_ _2400_ reg_data\[15\]\[31\] vssd1 vssd1
+ vccd1 vccd1 _2906_ sky130_fd_sc_hd__a32o_1
X_6272_ reg_data\[18\]\[30\] _1039_ _1063_ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__and3_1
X_9060_ clknet_leaf_63_i_clk _0204_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8011_ i_data[23] vssd1 vssd1 vccd1 vccd1 _3907_ sky130_fd_sc_hd__buf_2
X_5223_ reg_data\[4\]\[12\] _1824_ _1180_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__and3_1
X_5154_ reg_data\[27\]\[11\] _1199_ _1755_ _1756_ _1757_ vssd1 vssd1 vccd1 vccd1 _1758_
+ sky130_fd_sc_hd__a2111o_1
X_5085_ reg_data\[0\]\[10\] _1174_ _1688_ _1689_ _1690_ vssd1 vssd1 vccd1 vccd1 _1691_
+ sky130_fd_sc_hd__a2111o_1
X_8913_ clknet_leaf_21_i_clk _0057_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_9893_ clknet_leaf_75_i_clk _0963_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_8844_ reg_data\[11\]\[26\] i_data[26] _4346_ vssd1 vssd1 vccd1 vccd1 _4353_ sky130_fd_sc_hd__mux2_1
X_8775_ _4316_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__clkbuf_1
X_5987_ _2550_ _2554_ _2559_ _2564_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__or4_1
X_7726_ _3744_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__clkbuf_1
X_4938_ reg_data\[14\]\[8\] _1253_ _1379_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__and3_1
X_7657_ _3260_ reg_data\[24\]\[28\] _3699_ vssd1 vssd1 vccd1 vccd1 _3708_ sky130_fd_sc_hd__mux2_1
X_4869_ reg_data\[25\]\[7\] _1037_ _1478_ _1479_ _1481_ vssd1 vssd1 vccd1 vccd1 _1482_
+ sky130_fd_sc_hd__a2111o_1
X_6608_ _3110_ vssd1 vssd1 vccd1 vccd1 o_data2[24] sky130_fd_sc_hd__buf_2
X_7588_ reg_data\[23\]\[28\] _3187_ _3662_ vssd1 vssd1 vccd1 vccd1 _3671_ sky130_fd_sc_hd__mux2_1
X_9327_ clknet_leaf_30_i_clk _0471_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6539_ _3073_ vssd1 vssd1 vccd1 vccd1 o_data1[24] sky130_fd_sc_hd__buf_2
X_9258_ clknet_leaf_56_i_clk _0402_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_9189_ clknet_leaf_63_i_clk _0333_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8209_ _4016_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__clkbuf_1
X_5910_ reg_data\[17\]\[23\] _2489_ _1395_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__and3_1
X_6890_ _3297_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__clkbuf_1
X_5841_ reg_data\[18\]\[22\] _2422_ _2120_ vssd1 vssd1 vccd1 vccd1 _2423_ sky130_fd_sc_hd__and3_1
X_5772_ reg_data\[13\]\[21\] _2183_ _2299_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__and3_1
X_8560_ reg_data\[1\]\[20\] _3170_ _4202_ vssd1 vssd1 vccd1 vccd1 _4203_ sky130_fd_sc_hd__mux2_1
X_7511_ _3252_ reg_data\[21\]\[24\] _3625_ vssd1 vssd1 vccd1 vccd1 _3630_ sky130_fd_sc_hd__mux2_1
X_8491_ _4143_ vssd1 vssd1 vccd1 vccd1 _4166_ sky130_fd_sc_hd__clkbuf_8
X_4723_ reg_data\[18\]\[4\] _1159_ _1168_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__and3_1
X_7442_ _3592_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__clkbuf_1
X_4654_ reg_data\[21\]\[3\] _1272_ _1273_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__and3_1
X_7373_ reg_data\[3\]\[24\] _3179_ _3551_ vssd1 vssd1 vccd1 vccd1 _3556_ sky130_fd_sc_hd__mux2_1
X_4585_ _0997_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__clkbuf_2
X_6324_ reg_data\[17\]\[31\] _1058_ _1238_ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__and3_1
X_9112_ clknet_leaf_13_i_clk _0256_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_9043_ clknet_leaf_33_i_clk _0187_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6255_ reg_data\[12\]\[29\] _2562_ _1289_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__and3_1
X_5206_ _1785_ _1796_ _1802_ _1808_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__or4_1
X_6186_ _2756_ vssd1 vssd1 vccd1 vccd1 rdata1\[28\] sky130_fd_sc_hd__clkbuf_1
X_5137_ reg_data\[18\]\[11\] _1159_ _1513_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__and3_1
X_5068_ reg_data\[8\]\[10\] _1116_ _1119_ reg_data\[10\]\[10\] _1674_ vssd1 vssd1
+ vccd1 vccd1 _1675_ sky130_fd_sc_hd__a221o_1
X_9876_ clknet_leaf_53_i_clk _0946_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8827_ reg_data\[11\]\[18\] i_data[18] _4335_ vssd1 vssd1 vccd1 vccd1 _4344_ sky130_fd_sc_hd__mux2_1
X_8758_ _4307_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__clkbuf_1
X_7709_ _3243_ reg_data\[25\]\[20\] _3735_ vssd1 vssd1 vccd1 vccd1 _3736_ sky130_fd_sc_hd__mux2_1
X_8689_ reg_data\[19\]\[17\] _3164_ _4263_ vssd1 vssd1 vccd1 vccd1 _4271_ sky130_fd_sc_hd__mux2_1
X_4370_ _1001_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__buf_4
X_6040_ reg_data\[7\]\[25\] _2433_ _2613_ _2614_ _2615_ vssd1 vssd1 vccd1 vccd1 _2616_
+ sky130_fd_sc_hd__a2111o_1
X_7991_ _3893_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__clkbuf_1
X_6942_ _3233_ reg_data\[10\]\[15\] _3320_ vssd1 vssd1 vccd1 vccd1 _3326_ sky130_fd_sc_hd__mux2_1
X_9730_ clknet_leaf_7_i_clk _0874_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6873_ _3288_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__clkbuf_1
X_9661_ clknet_leaf_3_i_clk _0805_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_5824_ reg_data\[16\]\[22\] _2405_ _2406_ reg_data\[9\]\[22\] vssd1 vssd1 vccd1 vccd1
+ _2407_ sky130_fd_sc_hd__a22o_1
X_8612_ _4230_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__clkbuf_1
X_9592_ clknet_leaf_69_i_clk _0736_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8543_ reg_data\[1\]\[12\] _3154_ _4191_ vssd1 vssd1 vccd1 vccd1 _4194_ sky130_fd_sc_hd__mux2_1
X_5755_ reg_data\[8\]\[21\] _1797_ _1798_ reg_data\[10\]\[21\] _2339_ vssd1 vssd1
+ vccd1 vccd1 _2340_ sky130_fd_sc_hd__a221o_1
X_5686_ reg_data\[13\]\[20\] _2214_ _2102_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__and3_1
X_8474_ _4157_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__clkbuf_1
X_4706_ reg_data\[7\]\[4\] _1081_ _1322_ _1323_ _1324_ vssd1 vssd1 vccd1 vccd1 _1325_
+ sky130_fd_sc_hd__a2111o_1
X_7425_ _3583_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__clkbuf_1
X_4637_ reg_data\[13\]\[3\] _1089_ _1257_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__and3_1
X_4568_ rs2_mux\[0\] _1006_ rs2_mux\[2\] rs2_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1190_
+ sky130_fd_sc_hd__and4_2
X_7356_ reg_data\[3\]\[16\] _3162_ _3540_ vssd1 vssd1 vccd1 vccd1 _3547_ sky130_fd_sc_hd__mux2_1
X_6307_ reg_data\[13\]\[30\] _1177_ _2299_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__and3_1
X_4499_ _1020_ _1035_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__and2_4
X_7287_ _3510_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__clkbuf_1
X_6238_ reg_data\[24\]\[29\] _2409_ _2410_ reg_data\[28\]\[29\] _2806_ vssd1 vssd1
+ vccd1 vccd1 _2807_ sky130_fd_sc_hd__a221o_1
X_9026_ clknet_leaf_62_i_clk _0170_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6169_ reg_data\[4\]\[28\] _2325_ _2469_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__and3_1
X_9859_ clknet_leaf_67_i_clk _0929_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_5_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5540_ reg_data\[7\]\[17\] _1827_ _2129_ _2130_ _2131_ vssd1 vssd1 vccd1 vccd1 _2132_
+ sky130_fd_sc_hd__a2111o_1
X_5471_ _0999_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__buf_2
X_7210_ _3469_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__clkbuf_1
X_4422_ reg_data\[21\]\[2\] _1042_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__and3_1
X_8190_ _4006_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__clkbuf_1
X_7141_ reg_data\[7\]\[11\] _3152_ _3431_ vssd1 vssd1 vccd1 vccd1 _3433_ sky130_fd_sc_hd__mux2_1
X_7072_ _3225_ reg_data\[8\]\[11\] _3394_ vssd1 vssd1 vccd1 vccd1 _3396_ sky130_fd_sc_hd__mux2_1
X_6023_ _2591_ _2595_ _2597_ _2599_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__or4_1
X_7974_ i_data[11] vssd1 vssd1 vccd1 vccd1 _3882_ sky130_fd_sc_hd__buf_2
X_9713_ clknet_leaf_35_i_clk _0857_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6925_ _3216_ reg_data\[10\]\[7\] _3309_ vssd1 vssd1 vccd1 vccd1 _3317_ sky130_fd_sc_hd__mux2_1
X_9644_ clknet_leaf_28_i_clk _0788_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6856_ _3279_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__clkbuf_1
X_5807_ reg_data\[7\]\[22\] _2386_ _2387_ _2388_ _2389_ vssd1 vssd1 vccd1 vccd1 _2390_
+ sky130_fd_sc_hd__a2111o_1
X_9575_ clknet_leaf_56_i_clk _0719_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6787_ _3234_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__clkbuf_1
X_5738_ _1047_ vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__clkbuf_4
X_8526_ reg_data\[1\]\[4\] _3137_ _4180_ vssd1 vssd1 vccd1 vccd1 _4185_ sky130_fd_sc_hd__mux2_1
X_5669_ _1047_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__clkbuf_4
X_8457_ _4148_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__clkbuf_1
X_7408_ _3574_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__clkbuf_1
X_8388_ _3865_ reg_data\[17\]\[3\] _4108_ vssd1 vssd1 vccd1 vccd1 _4112_ sky130_fd_sc_hd__mux2_1
X_7339_ reg_data\[3\]\[8\] _3145_ _3529_ vssd1 vssd1 vccd1 vccd1 _3538_ sky130_fd_sc_hd__mux2_1
X_9009_ clknet_leaf_21_i_clk _0153_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_4971_ _1566_ _1570_ _1574_ _1580_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__or4_1
X_6710_ _3180_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__clkbuf_1
X_7690_ _3225_ reg_data\[25\]\[11\] _3724_ vssd1 vssd1 vccd1 vccd1 _3726_ sky130_fd_sc_hd__mux2_1
X_6641_ reg_data\[4\]\[2\] _3133_ _3129_ vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__mux2_1
X_9360_ clknet_leaf_31_i_clk _0504_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_8311_ i_rd[4] _3121_ _3197_ vssd1 vssd1 vccd1 vccd1 _4070_ sky130_fd_sc_hd__and3_2
X_6572_ _3091_ vssd1 vssd1 vccd1 vccd1 o_data2[7] sky130_fd_sc_hd__buf_2
X_9291_ clknet_leaf_58_i_clk _0435_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5523_ reg_data\[22\]\[17\] _1679_ _1622_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__and3_1
X_8242_ _4033_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__clkbuf_1
X_5454_ reg_data\[1\]\[16\] _1729_ _1793_ _1794_ reg_data\[15\]\[16\] vssd1 vssd1
+ vccd1 vccd1 _2049_ sky130_fd_sc_hd__a32o_1
X_4405_ _0994_ _1027_ _1028_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__a31o_1
X_8173_ _3923_ reg_data\[13\]\[31\] _3962_ vssd1 vssd1 vccd1 vccd1 _3997_ sky130_fd_sc_hd__mux2_1
X_5385_ reg_data\[4\]\[15\] _1718_ _1863_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__and3_1
X_7124_ reg_data\[7\]\[3\] _3135_ _3420_ vssd1 vssd1 vccd1 vccd1 _3424_ sky130_fd_sc_hd__mux2_1
X_7055_ _3208_ reg_data\[8\]\[3\] _3383_ vssd1 vssd1 vccd1 vccd1 _3387_ sky130_fd_sc_hd__mux2_1
X_6006_ reg_data\[6\]\[25\] _2207_ _2323_ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__and3_1
X_7957_ _3870_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__clkbuf_1
X_6908_ _3121_ _3124_ _3306_ vssd1 vssd1 vccd1 vccd1 _3307_ sky130_fd_sc_hd__and3_2
X_7888_ _3218_ reg_data\[28\]\[8\] _3822_ vssd1 vssd1 vccd1 vccd1 _3831_ sky130_fd_sc_hd__mux2_1
X_6839_ _3268_ _3269_ vssd1 vssd1 vccd1 vccd1 _3270_ sky130_fd_sc_hd__nor2_4
X_9627_ clknet_leaf_7_i_clk _0771_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_9558_ clknet_leaf_16_i_clk _0702_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_9489_ clknet_leaf_21_i_clk _0633_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_8509_ _4175_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_70_i_clk clknet_3_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_23_i_clk clknet_3_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5170_ reg_data\[30\]\[12\] _1597_ _1254_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_38_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_8860_ clknet_leaf_4_i_clk _0004_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_7811_ _3210_ reg_data\[27\]\[4\] _3785_ vssd1 vssd1 vccd1 vccd1 _3790_ sky130_fd_sc_hd__mux2_1
X_8791_ _4325_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__clkbuf_1
X_7742_ _3753_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__clkbuf_1
X_4954_ reg_data\[17\]\[8\] _1272_ _1395_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__and3_1
X_4885_ reg_data\[23\]\[7\] _1099_ _1101_ reg_data\[19\]\[7\] vssd1 vssd1 vccd1 vccd1
+ _1498_ sky130_fd_sc_hd__a22o_1
X_9412_ clknet_leaf_62_i_clk _0556_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_7673_ _3208_ reg_data\[25\]\[3\] _3713_ vssd1 vssd1 vccd1 vccd1 _3717_ sky130_fd_sc_hd__mux2_1
X_6624_ i_rd[0] i_rd[1] i_rd[2] vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__or3_1
X_6555_ rs2\[1\] rs2\[3\] _3081_ vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__nand3_4
X_9343_ clknet_leaf_72_i_clk _0487_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5506_ reg_data\[0\]\[17\] _1775_ _2095_ _2096_ _2098_ vssd1 vssd1 vccd1 vccd1 _2099_
+ sky130_fd_sc_hd__a2111o_1
X_9274_ clknet_leaf_61_i_clk _0418_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8225_ _3907_ reg_data\[14\]\[23\] _4021_ vssd1 vssd1 vccd1 vccd1 _4025_ sky130_fd_sc_hd__mux2_1
X_6486_ rs1\[1\] rs1\[3\] _3044_ vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__nand3_4
X_5437_ reg_data\[25\]\[16\] _1764_ _2029_ _2030_ _2031_ vssd1 vssd1 vccd1 vccd1 _2032_
+ sky130_fd_sc_hd__a2111o_1
X_8156_ _3988_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__clkbuf_1
X_5368_ reg_data\[1\]\[14\] _1904_ _1905_ reg_data\[15\]\[14\] vssd1 vssd1 vccd1 vccd1
+ _1966_ sky130_fd_sc_hd__a22o_1
X_8087_ _3951_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__clkbuf_1
X_7107_ _3260_ reg_data\[8\]\[28\] _3405_ vssd1 vssd1 vccd1 vccd1 _3414_ sky130_fd_sc_hd__mux2_1
X_5299_ _1886_ _1890_ _1894_ _1898_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__or4_1
X_7038_ _3376_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__clkbuf_1
X_8989_ clknet_leaf_3_i_clk _0133_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_4670_ reg_data\[12\]\[3\] _1189_ _1289_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__and3_1
X_6340_ reg_data\[2\]\[31\] _1021_ _2396_ _2397_ reg_data\[11\]\[31\] vssd1 vssd1
+ vccd1 vccd1 _2905_ sky130_fd_sc_hd__a32o_1
X_6271_ reg_data\[25\]\[30\] _2370_ _2835_ _2836_ _2837_ vssd1 vssd1 vccd1 vccd1 _2838_
+ sky130_fd_sc_hd__a2111o_1
X_8010_ _3906_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__clkbuf_1
X_5222_ _1000_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__clkbuf_4
X_5153_ reg_data\[1\]\[11\] _1298_ _1299_ reg_data\[15\]\[11\] vssd1 vssd1 vccd1 vccd1
+ _1757_ sky130_fd_sc_hd__a22o_1
X_5084_ reg_data\[5\]\[10\] _1179_ _1285_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__and3_1
X_8912_ clknet_leaf_22_i_clk _0056_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_9892_ clknet_leaf_74_i_clk _0962_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8843_ _4352_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__clkbuf_1
X_8774_ _3911_ reg_data\[29\]\[25\] _4310_ vssd1 vssd1 vccd1 vccd1 _4316_ sky130_fd_sc_hd__mux2_1
X_5986_ reg_data\[7\]\[24\] _2433_ _2560_ _2561_ _2563_ vssd1 vssd1 vccd1 vccd1 _2564_
+ sky130_fd_sc_hd__a2111o_1
X_7725_ _3260_ reg_data\[25\]\[28\] _3735_ vssd1 vssd1 vccd1 vccd1 _3744_ sky130_fd_sc_hd__mux2_1
X_4937_ reg_data\[0\]\[8\] _1070_ _1545_ _1546_ _1547_ vssd1 vssd1 vccd1 vccd1 _1548_
+ sky130_fd_sc_hd__a2111o_1
X_7656_ _3707_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__clkbuf_1
X_4868_ reg_data\[17\]\[7\] _1480_ _1108_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__and3_1
X_6607_ r_data2\[24\] _3105_ vssd1 vssd1 vccd1 vccd1 _3110_ sky130_fd_sc_hd__and2_1
X_7587_ _3670_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__clkbuf_1
X_9326_ clknet_leaf_28_i_clk _0470_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_4799_ _1399_ _1405_ _1410_ _1414_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__or4_2
X_6538_ r_data1\[24\] _3068_ vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__and2_1
X_6469_ reg_data\[0\]\[1\] _1173_ _3026_ _3027_ _3028_ vssd1 vssd1 vccd1 vccd1 _3029_
+ sky130_fd_sc_hd__a2111o_1
X_9257_ clknet_leaf_60_i_clk _0401_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_9188_ clknet_leaf_63_i_clk _0332_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8208_ _3890_ reg_data\[14\]\[15\] _4010_ vssd1 vssd1 vccd1 vccd1 _4016_ sky130_fd_sc_hd__mux2_1
X_8139_ _3979_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__clkbuf_1
X_5840_ _1142_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__clkbuf_4
X_5771_ reg_data\[0\]\[21\] _1821_ _2352_ _2353_ _2354_ vssd1 vssd1 vccd1 vccd1 _2355_
+ sky130_fd_sc_hd__a2111o_1
X_7510_ _3629_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__clkbuf_1
X_8490_ _4165_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__clkbuf_1
X_4722_ reg_data\[25\]\[4\] _1141_ _1336_ _1337_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_
+ sky130_fd_sc_hd__a2111o_1
X_7441_ _3252_ reg_data\[20\]\[24\] _3587_ vssd1 vssd1 vccd1 vccd1 _3592_ sky130_fd_sc_hd__mux2_1
X_4653_ _1144_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__clkbuf_4
X_7372_ _3555_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__clkbuf_1
X_4584_ _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__buf_4
X_6323_ reg_data\[21\]\[31\] _2372_ _1043_ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__and3_1
X_9111_ clknet_leaf_14_i_clk _0255_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_9042_ clknet_leaf_32_i_clk _0186_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6254_ reg_data\[14\]\[29\] _2301_ _1344_ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__and3_1
X_5205_ reg_data\[24\]\[12\] _1803_ _1804_ reg_data\[28\]\[12\] _1807_ vssd1 vssd1
+ vccd1 vccd1 _1808_ sky130_fd_sc_hd__a221o_1
X_6185_ _2747_ _2751_ _2753_ _2755_ vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__or4_1
X_5136_ reg_data\[25\]\[11\] _1141_ _1737_ _1738_ _1739_ vssd1 vssd1 vccd1 vccd1 _1740_
+ sky130_fd_sc_hd__a2111o_1
X_5067_ reg_data\[16\]\[10\] _1121_ _1123_ reg_data\[9\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _1674_ sky130_fd_sc_hd__a22o_1
X_9875_ clknet_leaf_58_i_clk _0945_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_8826_ _4343_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__clkbuf_1
X_5969_ reg_data\[22\]\[24\] _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__and3_1
X_8757_ _3894_ reg_data\[29\]\[17\] _4299_ vssd1 vssd1 vccd1 vccd1 _4307_ sky130_fd_sc_hd__mux2_1
X_7708_ _3712_ vssd1 vssd1 vccd1 vccd1 _3735_ sky130_fd_sc_hd__buf_4
X_8688_ _4270_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__clkbuf_1
X_7639_ _3698_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__clkbuf_1
X_9309_ clknet_leaf_67_i_clk _0453_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_7990_ _3892_ reg_data\[9\]\[16\] _3880_ vssd1 vssd1 vccd1 vccd1 _3893_ sky130_fd_sc_hd__mux2_1
X_6941_ _3325_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__clkbuf_1
X_6872_ reg_data\[2\]\[15\] _3160_ _3282_ vssd1 vssd1 vccd1 vccd1 _3288_ sky130_fd_sc_hd__mux2_1
X_9660_ clknet_leaf_11_i_clk _0804_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_5823_ _1122_ vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__buf_2
X_9591_ clknet_leaf_42_i_clk _0735_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_8611_ _3884_ reg_data\[12\]\[12\] _4227_ vssd1 vssd1 vccd1 vccd1 _4230_ sky130_fd_sc_hd__mux2_1
X_8542_ _4193_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__clkbuf_1
X_5754_ reg_data\[16\]\[21\] _1799_ _1800_ reg_data\[9\]\[21\] vssd1 vssd1 vccd1 vccd1
+ _2339_ sky130_fd_sc_hd__a22o_1
X_5685_ reg_data\[12\]\[20\] _1986_ _2271_ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__and3_1
X_8473_ _3882_ reg_data\[18\]\[11\] _4155_ vssd1 vssd1 vccd1 vccd1 _4157_ sky130_fd_sc_hd__mux2_1
X_4705_ reg_data\[14\]\[4\] _1089_ _1090_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__and3_1
X_4636_ _1086_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__clkbuf_4
X_7424_ _3235_ reg_data\[20\]\[16\] _3576_ vssd1 vssd1 vccd1 vccd1 _3583_ sky130_fd_sc_hd__mux2_1
X_7355_ _3546_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_1
X_6306_ reg_data\[0\]\[30\] _2427_ _2869_ _2870_ _2871_ vssd1 vssd1 vccd1 vccd1 _2872_
+ sky130_fd_sc_hd__a2111o_1
X_4567_ _1171_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__clkbuf_2
X_4498_ _1120_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__clkbuf_4
X_7286_ reg_data\[5\]\[15\] _3160_ _3504_ vssd1 vssd1 vccd1 vccd1 _3510_ sky130_fd_sc_hd__mux2_1
X_6237_ reg_data\[26\]\[29\] _2411_ _2412_ reg_data\[29\]\[29\] vssd1 vssd1 vccd1
+ vccd1 _2806_ sky130_fd_sc_hd__a22o_1
X_9025_ clknet_leaf_73_i_clk _0169_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6168_ reg_data\[6\]\[28\] _2207_ _2323_ vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__and3_1
X_5119_ reg_data\[13\]\[11\] _1608_ _1257_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__and3_1
X_6099_ reg_data\[27\]\[26\] _2439_ _2670_ _2671_ _2672_ vssd1 vssd1 vccd1 vccd1 _2673_
+ sky130_fd_sc_hd__a2111o_1
X_9858_ clknet_leaf_69_i_clk _0928_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8809_ _4334_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__clkbuf_1
X_9789_ clknet_leaf_55_i_clk rdata1\[5\] vssd1 vssd1 vccd1 vccd1 r_data1\[5\] sky130_fd_sc_hd__dfxtp_1
X_5470_ reg_data\[6\]\[16\] _1951_ _1632_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__and3_1
X_4421_ _1043_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__buf_4
X_7140_ _3432_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
X_7071_ _3395_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
X_6022_ reg_data\[24\]\[25\] _2409_ _2410_ reg_data\[28\]\[25\] _2598_ vssd1 vssd1
+ vccd1 vccd1 _2599_ sky130_fd_sc_hd__a221o_1
X_7973_ _3881_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__clkbuf_1
X_9712_ clknet_leaf_35_i_clk _0856_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6924_ _3316_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__clkbuf_1
X_9643_ clknet_leaf_44_i_clk _0787_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6855_ reg_data\[2\]\[7\] _3143_ _3271_ vssd1 vssd1 vccd1 vccd1 _3279_ sky130_fd_sc_hd__mux2_1
X_5806_ reg_data\[13\]\[22\] _2214_ _2102_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__and3_1
X_9574_ clknet_leaf_55_i_clk _0718_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6786_ _3233_ reg_data\[22\]\[15\] _3223_ vssd1 vssd1 vccd1 vccd1 _3234_ sky130_fd_sc_hd__mux2_1
X_5737_ reg_data\[3\]\[21\] _1770_ _2319_ _2320_ _2321_ vssd1 vssd1 vccd1 vccd1 _2322_
+ sky130_fd_sc_hd__a2111o_1
X_8525_ _4184_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__clkbuf_1
X_8456_ _3865_ reg_data\[18\]\[3\] _4144_ vssd1 vssd1 vccd1 vccd1 _4148_ sky130_fd_sc_hd__mux2_1
X_7407_ _3218_ reg_data\[20\]\[8\] _3565_ vssd1 vssd1 vccd1 vccd1 _3574_ sky130_fd_sc_hd__mux2_1
X_5668_ _2255_ vssd1 vssd1 vccd1 vccd1 rdata2\[19\] sky130_fd_sc_hd__clkbuf_1
X_8387_ _4111_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__clkbuf_1
X_5599_ reg_data\[23\]\[18\] _1834_ _1835_ reg_data\[19\]\[18\] vssd1 vssd1 vccd1
+ vccd1 _2189_ sky130_fd_sc_hd__a22o_1
X_4619_ _1043_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__clkbuf_4
X_7338_ _3537_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__clkbuf_1
X_7269_ reg_data\[5\]\[7\] _3143_ _3493_ vssd1 vssd1 vccd1 vccd1 _3501_ sky130_fd_sc_hd__mux2_1
X_9008_ clknet_leaf_22_i_clk _0152_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_4970_ reg_data\[7\]\[8\] _1185_ _1577_ _1578_ _1579_ vssd1 vssd1 vccd1 vccd1 _1580_
+ sky130_fd_sc_hd__a2111o_1
X_6640_ i_data[2] vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__clkbuf_4
X_6571_ r_data2\[7\] _3083_ vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__and2_1
X_8310_ _4069_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__clkbuf_1
X_5522_ _2114_ vssd1 vssd1 vccd1 vccd1 rdata1\[17\] sky130_fd_sc_hd__clkbuf_1
X_9290_ clknet_leaf_54_i_clk _0434_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8241_ _3923_ reg_data\[14\]\[31\] _3998_ vssd1 vssd1 vccd1 vccd1 _4033_ sky130_fd_sc_hd__mux2_1
X_5453_ reg_data\[2\]\[16\] _1613_ _1790_ _1791_ reg_data\[11\]\[16\] vssd1 vssd1
+ vccd1 vccd1 _2048_ sky130_fd_sc_hd__a32o_1
X_4404_ i_rs_valid rs1\[2\] vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__nor2_1
X_8172_ _3996_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__clkbuf_1
X_5384_ reg_data\[6\]\[15\] _1600_ _1716_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__and3_1
X_7123_ _3423_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
X_7054_ _3386_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_1
X_6005_ reg_data\[3\]\[25\] _2376_ _2579_ _2580_ _2581_ vssd1 vssd1 vccd1 vccd1 _2582_
+ sky130_fd_sc_hd__a2111o_1
X_7956_ _3869_ reg_data\[9\]\[5\] _3859_ vssd1 vssd1 vccd1 vccd1 _3870_ sky130_fd_sc_hd__mux2_1
X_7887_ _3830_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__clkbuf_1
X_6907_ i_rd[4] _3122_ vssd1 vssd1 vccd1 vccd1 _3306_ sky130_fd_sc_hd__xor2_1
X_6838_ i_rd[4] _3196_ _3124_ vssd1 vssd1 vccd1 vccd1 _3269_ sky130_fd_sc_hd__or3_4
X_9626_ clknet_leaf_9_i_clk _0770_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_9557_ clknet_leaf_16_i_clk _0701_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_8508_ _3917_ reg_data\[18\]\[28\] _4166_ vssd1 vssd1 vccd1 vccd1 _4175_ sky130_fd_sc_hd__mux2_1
X_6769_ i_data[10] vssd1 vssd1 vccd1 vccd1 _3222_ sky130_fd_sc_hd__buf_2
X_9488_ clknet_leaf_22_i_clk _0632_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_8439_ _4138_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_4_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_7810_ _3789_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__clkbuf_1
X_8790_ reg_data\[11\]\[0\] i_data[0] _4324_ vssd1 vssd1 vccd1 vccd1 _4325_ sky130_fd_sc_hd__mux2_1
X_7741_ _3208_ reg_data\[26\]\[3\] _3749_ vssd1 vssd1 vccd1 vccd1 _3753_ sky130_fd_sc_hd__mux2_1
X_4953_ reg_data\[22\]\[8\] _1143_ _1270_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__and3_1
X_7672_ _3716_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__clkbuf_1
X_9411_ clknet_leaf_60_i_clk _0555_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6623_ i_data[0] vssd1 vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__buf_4
X_4884_ _1482_ _1487_ _1492_ _1496_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__or4_1
X_6554_ rs2\[0\] rs2\[4\] rs2\[2\] vssd1 vssd1 vccd1 vccd1 _3081_ sky130_fd_sc_hd__and3_1
X_9342_ clknet_leaf_71_i_clk _0486_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6485_ rs1\[0\] rs1\[4\] rs1\[2\] vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__and3_1
X_5505_ reg_data\[5\]\[17\] _2097_ _1925_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__and3_1
X_9273_ clknet_leaf_69_i_clk _0417_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8224_ _4024_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__clkbuf_1
X_5436_ reg_data\[21\]\[16\] _1480_ _1240_ vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__and3_1
X_8155_ _3905_ reg_data\[13\]\[22\] _3985_ vssd1 vssd1 vccd1 vccd1 _3988_ sky130_fd_sc_hd__mux2_1
X_5367_ reg_data\[2\]\[14\] _1837_ _1901_ _1902_ reg_data\[11\]\[14\] vssd1 vssd1
+ vccd1 vccd1 _1965_ sky130_fd_sc_hd__a32o_1
X_8086_ _3905_ reg_data\[30\]\[22\] _3948_ vssd1 vssd1 vccd1 vccd1 _3951_ sky130_fd_sc_hd__mux2_1
X_7106_ _3413_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__clkbuf_1
X_5298_ reg_data\[7\]\[13\] _1827_ _1895_ _1896_ _1897_ vssd1 vssd1 vccd1 vccd1 _1898_
+ sky130_fd_sc_hd__a2111o_1
X_7037_ reg_data\[0\]\[28\] _3187_ _3367_ vssd1 vssd1 vccd1 vccd1 _3376_ sky130_fd_sc_hd__mux2_1
X_8988_ clknet_leaf_5_i_clk _0132_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_7939_ _3307_ _3601_ vssd1 vssd1 vccd1 vccd1 _3858_ sky130_fd_sc_hd__nand2_4
X_9609_ clknet_leaf_52_i_clk _0753_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6270_ reg_data\[21\]\[30\] _1058_ _2087_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__and3_1
X_5221_ reg_data\[5\]\[12\] _1460_ _1273_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__and3_1
X_5152_ reg_data\[2\]\[11\] _1002_ _1295_ _1296_ reg_data\[11\]\[11\] vssd1 vssd1
+ vccd1 vccd1 _1756_ sky130_fd_sc_hd__a32o_1
X_5083_ reg_data\[4\]\[10\] _1460_ _1407_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__and3_1
X_8911_ clknet_leaf_30_i_clk _0055_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_9891_ clknet_leaf_73_i_clk _0961_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8842_ reg_data\[11\]\[25\] i_data[25] _4346_ vssd1 vssd1 vccd1 vccd1 _4352_ sky130_fd_sc_hd__mux2_1
X_8773_ _4315_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__clkbuf_1
X_7724_ _3743_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__clkbuf_1
X_5985_ reg_data\[12\]\[24\] _2562_ _2016_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__and3_1
X_4936_ reg_data\[5\]\[8\] _1490_ _1250_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__and3_1
X_7655_ _3258_ reg_data\[24\]\[27\] _3699_ vssd1 vssd1 vccd1 vccd1 _3707_ sky130_fd_sc_hd__mux2_1
X_4867_ _1034_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__clkbuf_4
X_7586_ reg_data\[23\]\[27\] _3185_ _3662_ vssd1 vssd1 vccd1 vccd1 _3670_ sky130_fd_sc_hd__mux2_1
X_6606_ _3109_ vssd1 vssd1 vccd1 vccd1 o_data2[23] sky130_fd_sc_hd__buf_2
X_9325_ clknet_leaf_28_i_clk _0469_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6537_ _3072_ vssd1 vssd1 vccd1 vccd1 o_data1[23] sky130_fd_sc_hd__buf_2
X_4798_ reg_data\[7\]\[5\] _1185_ _1411_ _1412_ _1413_ vssd1 vssd1 vccd1 vccd1 _1414_
+ sky130_fd_sc_hd__a2111o_1
X_6468_ reg_data\[5\]\[1\] _1189_ _1338_ vssd1 vssd1 vccd1 vccd1 _3028_ sky130_fd_sc_hd__and3_1
X_9256_ clknet_leaf_56_i_clk _0400_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6399_ reg_data\[8\]\[0\] _1115_ _1118_ reg_data\[10\]\[0\] _2961_ vssd1 vssd1 vccd1
+ vccd1 _2962_ sky130_fd_sc_hd__a221o_1
X_9187_ clknet_leaf_64_i_clk _0331_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8207_ _4015_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__clkbuf_1
X_5419_ reg_data\[14\]\[15\] _1693_ _1958_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__and3_1
X_8138_ _3888_ reg_data\[13\]\[14\] _3974_ vssd1 vssd1 vccd1 vccd1 _3979_ sky130_fd_sc_hd__mux2_1
X_8069_ _3888_ reg_data\[30\]\[14\] _3937_ vssd1 vssd1 vccd1 vccd1 _3942_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_22_i_clk clknet_3_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_37_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5770_ reg_data\[5\]\[21\] _1824_ _1954_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__and3_1
X_4721_ reg_data\[21\]\[4\] _1150_ _1338_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__and3_1
X_7440_ _3591_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__clkbuf_1
X_4652_ _1142_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__clkbuf_4
X_7371_ reg_data\[3\]\[23\] _3177_ _3551_ vssd1 vssd1 vccd1 vccd1 _3555_ sky130_fd_sc_hd__mux2_1
X_9110_ clknet_leaf_16_i_clk _0254_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_4583_ _1138_ _1183_ _1156_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__and3_4
X_6322_ reg_data\[22\]\[31\] _1097_ _1047_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__and3_1
X_9041_ clknet_leaf_33_i_clk _0185_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6253_ reg_data\[13\]\[29\] _1177_ _2299_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__and3_1
X_5204_ reg_data\[26\]\[12\] _1805_ _1806_ reg_data\[29\]\[12\] vssd1 vssd1 vccd1
+ vccd1 _1807_ sky130_fd_sc_hd__a22o_1
X_6184_ reg_data\[24\]\[28\] _2409_ _2410_ reg_data\[28\]\[28\] _2754_ vssd1 vssd1
+ vccd1 vccd1 _2755_ sky130_fd_sc_hd__a221o_1
X_5135_ reg_data\[17\]\[11\] _1509_ _1275_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__and3_1
X_5066_ reg_data\[27\]\[10\] _1096_ _1670_ _1671_ _1672_ vssd1 vssd1 vccd1 vccd1 _1673_
+ sky130_fd_sc_hd__a2111o_1
X_9874_ clknet_leaf_53_i_clk _0944_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_8825_ reg_data\[11\]\[17\] i_data[17] _4335_ vssd1 vssd1 vccd1 vccd1 _4343_ sky130_fd_sc_hd__mux2_1
X_5968_ _2546_ vssd1 vssd1 vccd1 vccd1 rdata1\[24\] sky130_fd_sc_hd__clkbuf_1
X_8756_ _4306_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__clkbuf_1
X_7707_ _3734_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__clkbuf_1
X_4919_ reg_data\[16\]\[7\] _1219_ _1221_ reg_data\[9\]\[7\] vssd1 vssd1 vccd1 vccd1
+ _1531_ sky130_fd_sc_hd__a22o_1
X_5899_ reg_data\[2\]\[23\] _2219_ _2396_ _2397_ reg_data\[11\]\[23\] vssd1 vssd1
+ vccd1 vccd1 _2480_ sky130_fd_sc_hd__a32o_1
X_8687_ reg_data\[19\]\[16\] _3162_ _4263_ vssd1 vssd1 vccd1 vccd1 _4270_ sky130_fd_sc_hd__mux2_1
X_7638_ _3241_ reg_data\[24\]\[19\] _3688_ vssd1 vssd1 vccd1 vccd1 _3698_ sky130_fd_sc_hd__mux2_1
X_7569_ reg_data\[23\]\[19\] _3168_ _3651_ vssd1 vssd1 vccd1 vccd1 _3661_ sky130_fd_sc_hd__mux2_1
X_9308_ clknet_leaf_7_i_clk _0452_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_9239_ clknet_leaf_25_i_clk _0383_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_1__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_6940_ _3231_ reg_data\[10\]\[14\] _3320_ vssd1 vssd1 vccd1 vccd1 _3325_ sky130_fd_sc_hd__mux2_1
X_6871_ _3287_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__clkbuf_1
X_5822_ _1120_ vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__buf_2
X_9590_ clknet_leaf_40_i_clk _0734_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_8610_ _4229_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__clkbuf_1
X_8541_ reg_data\[1\]\[11\] _3152_ _4191_ vssd1 vssd1 vccd1 vccd1 _4193_ sky130_fd_sc_hd__mux2_1
X_5753_ reg_data\[27\]\[21\] _1786_ _2334_ _2335_ _2337_ vssd1 vssd1 vccd1 vccd1 _2338_
+ sky130_fd_sc_hd__a2111o_1
X_4704_ reg_data\[12\]\[4\] _1085_ _1128_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__and3_1
X_5684_ _1083_ vssd1 vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__clkbuf_4
X_8472_ _4156_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__clkbuf_1
X_7423_ _3582_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__clkbuf_1
X_4635_ reg_data\[12\]\[3\] _1085_ _1128_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__and3_1
X_4566_ reg_data\[12\]\[2\] _1186_ _1187_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__and3_1
X_7354_ reg_data\[3\]\[15\] _3160_ _3540_ vssd1 vssd1 vccd1 vccd1 _3546_ sky130_fd_sc_hd__mux2_1
X_6305_ reg_data\[5\]\[30\] _2430_ _1338_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__and3_1
X_4497_ _1097_ _1068_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__and2_4
X_9024_ clknet_leaf_74_i_clk _0168_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7285_ _3509_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__clkbuf_1
X_6236_ reg_data\[8\]\[29\] _2403_ _2404_ reg_data\[10\]\[29\] _2804_ vssd1 vssd1
+ vccd1 vccd1 _2805_ sky130_fd_sc_hd__a221o_1
X_6167_ reg_data\[3\]\[28\] _2376_ _2735_ _2736_ _2737_ vssd1 vssd1 vccd1 vccd1 _2738_
+ sky130_fd_sc_hd__a2111o_1
X_5118_ reg_data\[12\]\[11\] _1381_ _1606_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__and3_1
X_6098_ reg_data\[1\]\[26\] _2510_ _2511_ reg_data\[15\]\[26\] vssd1 vssd1 vccd1 vccd1
+ _2672_ sky130_fd_sc_hd__a22o_1
X_5049_ _1038_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__buf_2
X_9857_ clknet_leaf_67_i_clk rs2_mux\[4\] vssd1 vssd1 vccd1 vccd1 rs2\[4\] sky130_fd_sc_hd__dfxtp_1
X_8808_ reg_data\[11\]\[9\] i_data[9] _4324_ vssd1 vssd1 vccd1 vccd1 _4334_ sky130_fd_sc_hd__mux2_1
X_9788_ clknet_leaf_74_i_clk rdata1\[4\] vssd1 vssd1 vccd1 vccd1 r_data1\[4\] sky130_fd_sc_hd__dfxtp_2
X_8739_ _4297_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__clkbuf_1
X_4420_ rs1_mux\[0\] _1026_ rs1_mux\[2\] _1033_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__and4_4
X_7070_ _3222_ reg_data\[8\]\[10\] _3394_ vssd1 vssd1 vccd1 vccd1 _3395_ sky130_fd_sc_hd__mux2_1
X_6021_ reg_data\[26\]\[25\] _2411_ _2412_ reg_data\[29\]\[25\] vssd1 vssd1 vccd1
+ vccd1 _2598_ sky130_fd_sc_hd__a22o_1
X_7972_ _3879_ reg_data\[9\]\[10\] _3880_ vssd1 vssd1 vccd1 vccd1 _3881_ sky130_fd_sc_hd__mux2_1
X_9711_ clknet_leaf_36_i_clk _0855_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6923_ _3214_ reg_data\[10\]\[6\] _3309_ vssd1 vssd1 vccd1 vccd1 _3316_ sky130_fd_sc_hd__mux2_1
X_9642_ clknet_leaf_40_i_clk _0786_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6854_ _3278_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__clkbuf_1
X_5805_ reg_data\[12\]\[22\] _1986_ _2271_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__and3_1
X_6785_ i_data[15] vssd1 vssd1 vccd1 vccd1 _3233_ sky130_fd_sc_hd__buf_2
X_9573_ clknet_leaf_58_i_clk _0717_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5736_ reg_data\[30\]\[21\] _2204_ _1254_ vssd1 vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__and3_1
X_8524_ reg_data\[1\]\[3\] _3135_ _4180_ vssd1 vssd1 vccd1 vccd1 _4184_ sky130_fd_sc_hd__mux2_1
X_5667_ _2246_ _2250_ _2252_ _2254_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__or4_1
X_8455_ _4147_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__clkbuf_1
X_7406_ _3573_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__clkbuf_1
X_4618_ reg_data\[17\]\[3\] _1042_ _1238_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__and3_1
X_5598_ _2174_ _2178_ _2182_ _2187_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__or4_2
X_8386_ _3863_ reg_data\[17\]\[2\] _4108_ vssd1 vssd1 vccd1 vccd1 _4111_ sky130_fd_sc_hd__mux2_1
X_4549_ _0999_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__buf_2
X_7337_ reg_data\[3\]\[7\] _3143_ _3529_ vssd1 vssd1 vccd1 vccd1 _3537_ sky130_fd_sc_hd__mux2_1
X_7268_ _3500_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__clkbuf_1
X_9007_ clknet_leaf_29_i_clk _0151_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6219_ reg_data\[20\]\[29\] _2524_ _1059_ vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__and3_1
X_7199_ _3463_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__clkbuf_1
X_9909_ clknet_leaf_59_i_clk _0979_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6570_ _3090_ vssd1 vssd1 vccd1 vccd1 o_data2[6] sky130_fd_sc_hd__buf_2
X_5521_ _2105_ _2109_ _2111_ _2113_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__or4_1
X_8240_ _4032_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__clkbuf_1
X_5452_ reg_data\[23\]\[16\] _1787_ _1788_ reg_data\[19\]\[16\] vssd1 vssd1 vccd1
+ vccd1 _2047_ sky130_fd_sc_hd__a22o_1
X_4403_ i_rs1[0] i_rs1[1] i_rs1[2] vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__o21ai_1
X_8171_ _3921_ reg_data\[13\]\[30\] _3962_ vssd1 vssd1 vccd1 vccd1 _3996_ sky130_fd_sc_hd__mux2_1
X_5383_ reg_data\[3\]\[15\] _1770_ _1977_ _1978_ _1979_ vssd1 vssd1 vccd1 vccd1 _1980_
+ sky130_fd_sc_hd__a2111o_1
X_7122_ reg_data\[7\]\[2\] _3133_ _3420_ vssd1 vssd1 vccd1 vccd1 _3423_ sky130_fd_sc_hd__mux2_1
X_7053_ _3206_ reg_data\[8\]\[2\] _3383_ vssd1 vssd1 vccd1 vccd1 _3386_ sky130_fd_sc_hd__mux2_1
X_6004_ reg_data\[20\]\[25\] _2204_ _2035_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__and3_1
X_7955_ i_data[5] vssd1 vssd1 vccd1 vccd1 _3869_ sky130_fd_sc_hd__clkbuf_4
X_6906_ _3305_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__clkbuf_1
X_7886_ _3216_ reg_data\[28\]\[7\] _3822_ vssd1 vssd1 vccd1 vccd1 _3830_ sky130_fd_sc_hd__mux2_1
X_6837_ i_rd[0] i_rd[1] i_write i_reset_n vssd1 vssd1 vccd1 vccd1 _3268_ sky130_fd_sc_hd__nand4_4
X_9625_ clknet_leaf_9_i_clk _0769_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_9556_ clknet_leaf_16_i_clk _0700_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_8507_ _4174_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__clkbuf_1
X_6768_ _3221_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__clkbuf_1
X_9487_ clknet_leaf_30_i_clk _0631_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_5719_ _2290_ _2294_ _2298_ _2304_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__or4_2
X_6699_ i_data[21] vssd1 vssd1 vccd1 vccd1 _3173_ sky130_fd_sc_hd__clkbuf_4
X_8438_ _3915_ reg_data\[17\]\[27\] _4130_ vssd1 vssd1 vccd1 vccd1 _4138_ sky130_fd_sc_hd__mux2_1
X_8369_ _4101_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__clkbuf_1
X_4952_ _1562_ vssd1 vssd1 vccd1 vccd1 rdata1\[8\] sky130_fd_sc_hd__clkbuf_1
X_7740_ _3752_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__clkbuf_1
X_4883_ reg_data\[7\]\[7\] _1081_ _1493_ _1494_ _1495_ vssd1 vssd1 vccd1 vccd1 _1496_
+ sky130_fd_sc_hd__a2111o_1
X_7671_ _3206_ reg_data\[25\]\[2\] _3713_ vssd1 vssd1 vccd1 vccd1 _3716_ sky130_fd_sc_hd__mux2_1
X_6622_ _3117_ vssd1 vssd1 vccd1 vccd1 o_data2[31] sky130_fd_sc_hd__buf_2
X_9410_ clknet_leaf_59_i_clk _0554_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6553_ _3080_ vssd1 vssd1 vccd1 vccd1 o_data1[31] sky130_fd_sc_hd__buf_2
X_9341_ clknet_leaf_69_i_clk _0485_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_5504_ _1067_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__clkbuf_4
X_9272_ clknet_leaf_61_i_clk _0416_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6484_ _3043_ vssd1 vssd1 vccd1 vccd1 rdata2\[1\] sky130_fd_sc_hd__clkbuf_1
X_8223_ _3905_ reg_data\[14\]\[22\] _4021_ vssd1 vssd1 vccd1 vccd1 _4024_ sky130_fd_sc_hd__mux2_1
X_5435_ reg_data\[17\]\[16\] _1766_ _1708_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__and3_1
X_8154_ _3987_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__clkbuf_1
X_5366_ reg_data\[23\]\[14\] _1834_ _1835_ reg_data\[19\]\[14\] vssd1 vssd1 vccd1
+ vccd1 _1964_ sky130_fd_sc_hd__a22o_1
X_7105_ _3258_ reg_data\[8\]\[27\] _3405_ vssd1 vssd1 vccd1 vccd1 _3413_ sky130_fd_sc_hd__mux2_1
X_8085_ _3950_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__clkbuf_1
X_5297_ reg_data\[12\]\[13\] _1354_ _1226_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__and3_1
X_7036_ _3375_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__clkbuf_1
X_8987_ clknet_leaf_0_i_clk _0131_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_7938_ i_data[0] vssd1 vssd1 vccd1 vccd1 _3857_ sky130_fd_sc_hd__clkbuf_4
X_7869_ _3121_ _3197_ _3306_ vssd1 vssd1 vccd1 vccd1 _3820_ sky130_fd_sc_hd__or3_1
X_9608_ clknet_leaf_53_i_clk _0752_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_9539_ clknet_leaf_8_i_clk _0683_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_5220_ reg_data\[6\]\[12\] _1347_ _1632_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__and3_1
X_5151_ reg_data\[23\]\[11\] _1206_ _1209_ reg_data\[19\]\[11\] vssd1 vssd1 vccd1
+ vccd1 _1755_ sky130_fd_sc_hd__a22o_1
X_5082_ reg_data\[6\]\[10\] _1347_ _1632_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__and3_1
X_8910_ clknet_leaf_32_i_clk _0054_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_9890_ clknet_leaf_73_i_clk _0960_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8841_ _4351_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__clkbuf_1
X_8772_ _3909_ reg_data\[29\]\[24\] _4310_ vssd1 vssd1 vccd1 vccd1 _4315_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_3_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_7723_ _3258_ reg_data\[25\]\[27\] _3735_ vssd1 vssd1 vccd1 vccd1 _3743_ sky130_fd_sc_hd__mux2_1
X_5984_ _1000_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__buf_2
X_4935_ reg_data\[4\]\[8\] _1074_ _1248_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__and3_1
X_7654_ _3706_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__clkbuf_1
X_4866_ reg_data\[21\]\[7\] _1042_ _1044_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__and3_1
X_7585_ _3669_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__clkbuf_1
X_6605_ r_data2\[23\] _3105_ vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__and2_1
X_4797_ reg_data\[12\]\[5\] _1354_ _1226_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__and3_1
X_9324_ clknet_leaf_28_i_clk _0468_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6536_ r_data1\[23\] _3068_ vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__and2_1
X_6467_ reg_data\[4\]\[1\] _1175_ _1342_ vssd1 vssd1 vccd1 vccd1 _3027_ sky130_fd_sc_hd__and3_1
X_9255_ clknet_leaf_56_i_clk _0399_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6398_ reg_data\[16\]\[0\] _1120_ _1122_ reg_data\[9\]\[0\] vssd1 vssd1 vccd1 vccd1
+ _2961_ sky130_fd_sc_hd__a22o_1
X_9186_ clknet_leaf_66_i_clk _0330_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8206_ _3888_ reg_data\[14\]\[14\] _4010_ vssd1 vssd1 vccd1 vccd1 _4015_ sky130_fd_sc_hd__mux2_1
X_5418_ reg_data\[13\]\[15\] _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__and3_1
X_5349_ reg_data\[18\]\[14\] _1816_ _1513_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__and3_1
X_8137_ _3978_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__clkbuf_1
X_8068_ _3941_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__clkbuf_1
X_7019_ _3366_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__clkbuf_1
X_4720_ _1144_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__buf_2
X_4651_ reg_data\[22\]\[3\] _1143_ _1270_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__and3_1
X_7370_ _3554_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__clkbuf_1
X_4582_ reg_data\[1\]\[2\] _1202_ _1203_ reg_data\[15\]\[2\] vssd1 vssd1 vccd1 vccd1
+ _1204_ sky130_fd_sc_hd__a22o_1
X_6321_ _2886_ vssd1 vssd1 vccd1 vccd1 rdata2\[30\] sky130_fd_sc_hd__clkbuf_1
X_9040_ clknet_leaf_33_i_clk _0184_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6252_ reg_data\[0\]\[29\] _2427_ _2817_ _2818_ _2819_ vssd1 vssd1 vccd1 vccd1 _2820_
+ sky130_fd_sc_hd__a2111o_1
X_6183_ reg_data\[26\]\[28\] _2411_ _2412_ reg_data\[29\]\[28\] vssd1 vssd1 vccd1
+ vccd1 _2754_ sky130_fd_sc_hd__a22o_1
X_5203_ _1133_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__clkbuf_4
X_5134_ reg_data\[21\]\[11\] _1272_ _1273_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__and3_1
X_5065_ reg_data\[1\]\[10\] _1022_ _1109_ _1111_ reg_data\[15\]\[10\] vssd1 vssd1
+ vccd1 vccd1 _1672_ sky130_fd_sc_hd__a32o_1
X_9873_ clknet_leaf_58_i_clk _0943_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8824_ _4342_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__clkbuf_1
X_5967_ _2537_ _2541_ _2543_ _2545_ vssd1 vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__or4_1
X_8755_ _3892_ reg_data\[29\]\[16\] _4299_ vssd1 vssd1 vccd1 vccd1 _4306_ sky130_fd_sc_hd__mux2_1
X_7706_ _3241_ reg_data\[25\]\[19\] _3724_ vssd1 vssd1 vccd1 vccd1 _3734_ sky130_fd_sc_hd__mux2_1
X_8686_ _4269_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__clkbuf_1
X_4918_ reg_data\[27\]\[7\] _1199_ _1527_ _1528_ _1529_ vssd1 vssd1 vccd1 vccd1 _1530_
+ sky130_fd_sc_hd__a2111o_1
X_5898_ reg_data\[23\]\[23\] _2393_ _2394_ reg_data\[19\]\[23\] vssd1 vssd1 vccd1
+ vccd1 _2479_ sky130_fd_sc_hd__a22o_1
X_7637_ _3697_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__clkbuf_1
X_4849_ reg_data\[0\]\[6\] _1174_ _1459_ _1461_ _1462_ vssd1 vssd1 vccd1 vccd1 _1463_
+ sky130_fd_sc_hd__a2111o_1
X_7568_ _3660_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__clkbuf_1
X_7499_ _3623_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__clkbuf_1
X_6519_ r_data1\[15\] _3057_ vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__and2_1
X_9307_ clknet_leaf_67_i_clk _0451_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_9238_ clknet_leaf_23_i_clk _0382_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_9169_ clknet_leaf_21_i_clk _0313_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6870_ reg_data\[2\]\[14\] _3158_ _3282_ vssd1 vssd1 vccd1 vccd1 _3287_ sky130_fd_sc_hd__mux2_1
X_5821_ _1118_ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__buf_2
X_5752_ reg_data\[1\]\[21\] _2336_ _1793_ _1794_ reg_data\[15\]\[21\] vssd1 vssd1
+ vccd1 vccd1 _2337_ sky130_fd_sc_hd__a32o_1
X_8540_ _4192_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__clkbuf_1
X_4703_ reg_data\[13\]\[4\] _1253_ _1087_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__and3_1
X_5683_ reg_data\[14\]\[20\] _1867_ _2156_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__and3_1
X_8471_ _3879_ reg_data\[18\]\[10\] _4155_ vssd1 vssd1 vccd1 vccd1 _4156_ sky130_fd_sc_hd__mux2_1
X_7422_ _3233_ reg_data\[20\]\[15\] _3576_ vssd1 vssd1 vccd1 vccd1 _3582_ sky130_fd_sc_hd__mux2_1
X_4634_ reg_data\[14\]\[3\] _1253_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__and3_1
X_4565_ _0993_ _1006_ rs2_mux\[2\] rs2_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__and4_4
X_7353_ _3545_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__clkbuf_1
X_6304_ reg_data\[4\]\[30\] _1175_ _1342_ vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_21_i_clk clknet_3_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_9023_ clknet_leaf_73_i_clk _0167_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_4496_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__clkbuf_4
X_7284_ reg_data\[5\]\[14\] _3158_ _3504_ vssd1 vssd1 vccd1 vccd1 _3509_ sky130_fd_sc_hd__mux2_1
X_6235_ reg_data\[16\]\[29\] _2405_ _2406_ reg_data\[9\]\[29\] vssd1 vssd1 vccd1 vccd1
+ _2804_ sky130_fd_sc_hd__a22o_1
X_6166_ reg_data\[20\]\[28\] _2204_ _2035_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__and3_1
X_6097_ reg_data\[2\]\[26\] _2443_ _2507_ _2508_ reg_data\[11\]\[26\] vssd1 vssd1
+ vccd1 vccd1 _2671_ sky130_fd_sc_hd__a32o_1
X_5117_ reg_data\[14\]\[11\] _1253_ _1379_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_36_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5048_ reg_data\[25\]\[10\] _1037_ _1652_ _1653_ _1654_ vssd1 vssd1 vccd1 vccd1 _1655_
+ sky130_fd_sc_hd__a2111o_1
X_9856_ clknet_leaf_24_i_clk rs2_mux\[3\] vssd1 vssd1 vccd1 vccd1 rs2\[3\] sky130_fd_sc_hd__dfxtp_1
X_9787_ clknet_leaf_71_i_clk rdata1\[3\] vssd1 vssd1 vccd1 vccd1 r_data1\[3\] sky130_fd_sc_hd__dfxtp_1
X_8807_ _4333_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__clkbuf_1
X_6999_ _3344_ vssd1 vssd1 vccd1 vccd1 _3356_ sky130_fd_sc_hd__buf_6
X_8738_ _3875_ reg_data\[29\]\[8\] _4288_ vssd1 vssd1 vccd1 vccd1 _4297_ sky130_fd_sc_hd__mux2_1
X_8669_ _4260_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__clkbuf_1
X_6020_ reg_data\[8\]\[25\] _2403_ _2404_ reg_data\[10\]\[25\] _2596_ vssd1 vssd1
+ vccd1 vccd1 _2597_ sky130_fd_sc_hd__a221o_1
X_7971_ _3858_ vssd1 vssd1 vccd1 vccd1 _3880_ sky130_fd_sc_hd__buf_4
X_9710_ clknet_leaf_39_i_clk _0854_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6922_ _3315_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__clkbuf_1
X_9641_ clknet_leaf_41_i_clk _0785_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6853_ reg_data\[2\]\[6\] _3141_ _3271_ vssd1 vssd1 vccd1 vccd1 _3278_ sky130_fd_sc_hd__mux2_1
X_5804_ reg_data\[14\]\[22\] _1867_ _2156_ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__and3_1
X_9572_ clknet_leaf_60_i_clk _0716_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_6784_ _3232_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__clkbuf_1
X_5735_ reg_data\[20\]\[21\] _1918_ _1060_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__and3_1
X_8523_ _4183_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__clkbuf_1
X_8454_ _3863_ reg_data\[18\]\[2\] _4144_ vssd1 vssd1 vccd1 vccd1 _4147_ sky130_fd_sc_hd__mux2_1
X_5666_ reg_data\[24\]\[19\] _1847_ _1848_ reg_data\[28\]\[19\] _2253_ vssd1 vssd1
+ vccd1 vccd1 _2254_ sky130_fd_sc_hd__a221o_1
X_4617_ _1040_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__buf_4
X_7405_ _3216_ reg_data\[20\]\[7\] _3565_ vssd1 vssd1 vccd1 vccd1 _3573_ sky130_fd_sc_hd__mux2_1
X_5597_ reg_data\[7\]\[18\] _1827_ _2184_ _2185_ _2186_ vssd1 vssd1 vccd1 vccd1 _2187_
+ sky130_fd_sc_hd__a2111o_1
X_8385_ _4110_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__clkbuf_1
X_7336_ _3536_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__clkbuf_1
X_4548_ reg_data\[3\]\[2\] _1158_ _1161_ _1165_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_
+ sky130_fd_sc_hd__a2111o_1
X_4479_ reg_data\[23\]\[2\] _1099_ _1101_ reg_data\[19\]\[2\] vssd1 vssd1 vccd1 vccd1
+ _1102_ sky130_fd_sc_hd__a22o_1
X_7267_ reg_data\[5\]\[6\] _3141_ _3493_ vssd1 vssd1 vccd1 vccd1 _3500_ sky130_fd_sc_hd__mux2_1
X_6218_ reg_data\[18\]\[29\] _2261_ _1063_ vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__and3_1
X_9006_ clknet_leaf_29_i_clk _0150_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_7198_ reg_data\[6\]\[6\] _3141_ _3456_ vssd1 vssd1 vccd1 vccd1 _3463_ sky130_fd_sc_hd__mux2_1
X_6149_ _2708_ _2712_ _2716_ _2720_ vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__or4_4
X_9908_ clknet_leaf_56_i_clk _0978_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_9839_ clknet_leaf_36_i_clk rdata2\[23\] vssd1 vssd1 vccd1 vccd1 r_data2\[23\] sky130_fd_sc_hd__dfxtp_1
X_5520_ reg_data\[24\]\[17\] _1803_ _1804_ reg_data\[28\]\[17\] _2112_ vssd1 vssd1
+ vccd1 vccd1 _2113_ sky130_fd_sc_hd__a221o_1
X_5451_ _2032_ _2037_ _2041_ _2045_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__or4_1
X_4402_ i_rs1[0] i_rs1[2] i_rs1[1] vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__or3_1
X_8170_ _3995_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__clkbuf_1
X_5382_ reg_data\[20\]\[15\] _1597_ _1315_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__and3_1
X_7121_ _3422_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
X_7052_ _3385_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_1
X_6003_ reg_data\[30\]\[25\] _2524_ _1919_ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__and3_1
X_7954_ _3868_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__clkbuf_1
X_6905_ reg_data\[2\]\[31\] _3193_ _3270_ vssd1 vssd1 vccd1 vccd1 _3305_ sky130_fd_sc_hd__mux2_1
X_7885_ _3829_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__clkbuf_1
X_6836_ _3267_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__clkbuf_1
X_9624_ clknet_leaf_9_i_clk _0768_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_9555_ clknet_leaf_17_i_clk _0699_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6767_ _3220_ reg_data\[22\]\[9\] _3202_ vssd1 vssd1 vccd1 vccd1 _3221_ sky130_fd_sc_hd__mux2_1
X_8506_ _3915_ reg_data\[18\]\[27\] _4166_ vssd1 vssd1 vccd1 vccd1 _4174_ sky130_fd_sc_hd__mux2_1
X_5718_ reg_data\[7\]\[20\] _1827_ _2300_ _2302_ _2303_ vssd1 vssd1 vccd1 vccd1 _2304_
+ sky130_fd_sc_hd__a2111o_1
X_9486_ clknet_leaf_30_i_clk _0630_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6698_ _3172_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__clkbuf_1
X_8437_ _4137_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__clkbuf_1
X_5649_ _1151_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__clkbuf_4
X_8368_ _3913_ reg_data\[16\]\[26\] _4094_ vssd1 vssd1 vccd1 vccd1 _4101_ sky130_fd_sc_hd__mux2_1
X_7319_ reg_data\[5\]\[31\] _3193_ _3492_ vssd1 vssd1 vccd1 vccd1 _3527_ sky130_fd_sc_hd__mux2_1
X_8299_ _3913_ reg_data\[15\]\[26\] _4057_ vssd1 vssd1 vccd1 vccd1 _4064_ sky130_fd_sc_hd__mux2_1
X_4951_ _1553_ _1557_ _1559_ _1561_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__or4_4
X_7670_ _3715_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__clkbuf_1
X_4882_ reg_data\[12\]\[7\] _1089_ _1128_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__and3_1
X_6621_ r_data2\[31\] _3082_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__and2_1
X_9340_ clknet_leaf_71_i_clk _0484_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6552_ r_data1\[31\] _3045_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__and2_1
X_9271_ clknet_leaf_39_i_clk _0415_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5503_ reg_data\[4\]\[17\] _1718_ _1863_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__and3_1
X_6483_ _3034_ _3038_ _3040_ _3042_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__or4_2
X_8222_ _4023_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__clkbuf_1
X_5434_ reg_data\[22\]\[16\] _1536_ _1651_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__and3_1
X_8153_ _3903_ reg_data\[13\]\[21\] _3985_ vssd1 vssd1 vccd1 vccd1 _3987_ sky130_fd_sc_hd__mux2_1
X_7104_ _3412_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__clkbuf_1
X_5365_ _1946_ _1950_ _1956_ _1962_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__or4_1
X_8084_ _3903_ reg_data\[30\]\[21\] _3948_ vssd1 vssd1 vccd1 vccd1 _3950_ sky130_fd_sc_hd__mux2_1
X_5296_ reg_data\[14\]\[13\] _1693_ _1193_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__and3_1
X_7035_ reg_data\[0\]\[27\] _3185_ _3367_ vssd1 vssd1 vccd1 vccd1 _3375_ sky130_fd_sc_hd__mux2_1
X_8986_ clknet_leaf_12_i_clk _0130_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_7937_ _3856_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__clkbuf_1
X_7868_ _3819_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__clkbuf_1
X_6819_ i_data[26] vssd1 vssd1 vccd1 vccd1 _3256_ sky130_fd_sc_hd__buf_2
X_9607_ clknet_leaf_51_i_clk _0751_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_7799_ _3266_ reg_data\[26\]\[31\] _3748_ vssd1 vssd1 vccd1 vccd1 _3783_ sky130_fd_sc_hd__mux2_1
X_9538_ clknet_leaf_65_i_clk _0682_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_9469_ clknet_leaf_4_i_clk _0613_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_5150_ _1740_ _1745_ _1749_ _1753_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__or4_1
X_5081_ reg_data\[3\]\[10\] _1158_ _1684_ _1685_ _1686_ vssd1 vssd1 vccd1 vccd1 _1687_
+ sky130_fd_sc_hd__a2111o_1
X_8840_ reg_data\[11\]\[24\] i_data[24] _4346_ vssd1 vssd1 vccd1 vccd1 _4351_ sky130_fd_sc_hd__mux2_1
X_8771_ _4314_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__clkbuf_1
X_5983_ reg_data\[14\]\[24\] _2301_ _1958_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__and3_1
X_7722_ _3742_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__clkbuf_1
X_4934_ reg_data\[6\]\[8\] _1072_ _1048_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__and3_1
X_7653_ _3256_ reg_data\[24\]\[26\] _3699_ vssd1 vssd1 vccd1 vccd1 _3706_ sky130_fd_sc_hd__mux2_1
X_4865_ reg_data\[22\]\[7\] _1039_ _1236_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__and3_1
X_7584_ reg_data\[23\]\[26\] _3183_ _3662_ vssd1 vssd1 vccd1 vccd1 _3669_ sky130_fd_sc_hd__mux2_1
X_6604_ _3108_ vssd1 vssd1 vccd1 vccd1 o_data2[22] sky130_fd_sc_hd__buf_2
X_4796_ reg_data\[14\]\[5\] _1189_ _1193_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__and3_1
X_9323_ clknet_leaf_44_i_clk _0467_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6535_ _3071_ vssd1 vssd1 vccd1 vccd1 o_data1[22] sky130_fd_sc_hd__buf_2
X_9254_ clknet_leaf_55_i_clk _0398_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6466_ reg_data\[6\]\[1\] _2555_ _1270_ vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__and3_1
X_8205_ _4014_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__clkbuf_1
X_6397_ reg_data\[27\]\[0\] _1095_ _2957_ _2958_ _2959_ vssd1 vssd1 vccd1 vccd1 _2960_
+ sky130_fd_sc_hd__a2111o_1
X_9185_ clknet_leaf_6_i_clk _0329_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5417_ reg_data\[0\]\[15\] _1821_ _2010_ _2011_ _2012_ vssd1 vssd1 vccd1 vccd1 _2013_
+ sky130_fd_sc_hd__a2111o_1
X_5348_ reg_data\[25\]\[14\] _1810_ _1942_ _1944_ _1945_ vssd1 vssd1 vccd1 vccd1 _1946_
+ sky130_fd_sc_hd__a2111o_1
X_8136_ _3886_ reg_data\[13\]\[13\] _3974_ vssd1 vssd1 vccd1 vccd1 _3978_ sky130_fd_sc_hd__mux2_1
X_8067_ _3886_ reg_data\[30\]\[13\] _3937_ vssd1 vssd1 vccd1 vccd1 _3941_ sky130_fd_sc_hd__mux2_1
X_7018_ reg_data\[0\]\[19\] _3168_ _3356_ vssd1 vssd1 vccd1 vccd1 _3366_ sky130_fd_sc_hd__mux2_1
X_5279_ reg_data\[24\]\[13\] _1803_ _1804_ reg_data\[28\]\[13\] _1879_ vssd1 vssd1
+ vccd1 vccd1 _1880_ sky130_fd_sc_hd__a221o_1
X_8969_ clknet_leaf_52_i_clk _0113_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_4650_ _1151_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__clkbuf_4
X_6320_ _2877_ _2881_ _2883_ _2885_ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__or4_1
X_4581_ _1000_ rs2_mux\[2\] rs2_mux\[3\] _1156_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__and4_4
X_6251_ reg_data\[5\]\[29\] _2430_ _1338_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__and3_1
X_6182_ reg_data\[8\]\[28\] _2403_ _2404_ reg_data\[10\]\[28\] _2752_ vssd1 vssd1
+ vccd1 vccd1 _2753_ sky130_fd_sc_hd__a221o_1
X_5202_ _1131_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__clkbuf_4
X_5133_ reg_data\[22\]\[11\] _1679_ _1622_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__and3_1
X_5064_ reg_data\[2\]\[10\] _1613_ _1104_ _1106_ reg_data\[11\]\[10\] vssd1 vssd1
+ vccd1 vccd1 _1671_ sky130_fd_sc_hd__a32o_1
X_9872_ clknet_leaf_53_i_clk _0942_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8823_ reg_data\[11\]\[16\] i_data[16] _4335_ vssd1 vssd1 vccd1 vccd1 _4342_ sky130_fd_sc_hd__mux2_1
X_5966_ reg_data\[24\]\[24\] _2409_ _2410_ reg_data\[28\]\[24\] _2544_ vssd1 vssd1
+ vccd1 vccd1 _2545_ sky130_fd_sc_hd__a221o_1
X_8754_ _4305_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__clkbuf_1
X_5897_ _2463_ _2467_ _2472_ _2477_ vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__or4_1
X_7705_ _3733_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__clkbuf_1
X_8685_ reg_data\[19\]\[15\] _3160_ _4263_ vssd1 vssd1 vccd1 vccd1 _4269_ sky130_fd_sc_hd__mux2_1
X_4917_ reg_data\[1\]\[7\] _1298_ _1299_ reg_data\[15\]\[7\] vssd1 vssd1 vccd1 vccd1
+ _1529_ sky130_fd_sc_hd__a22o_1
X_7636_ _3239_ reg_data\[24\]\[18\] _3688_ vssd1 vssd1 vccd1 vccd1 _3697_ sky130_fd_sc_hd__mux2_1
X_4848_ reg_data\[5\]\[6\] _1179_ _1285_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__and3_1
X_7567_ reg_data\[23\]\[18\] _3166_ _3651_ vssd1 vssd1 vccd1 vccd1 _3660_ sky130_fd_sc_hd__mux2_1
X_4779_ _1147_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__buf_4
X_9306_ clknet_leaf_9_i_clk _0450_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_7498_ _3239_ reg_data\[21\]\[18\] _3614_ vssd1 vssd1 vccd1 vccd1 _3623_ sky130_fd_sc_hd__mux2_1
X_6518_ _3062_ vssd1 vssd1 vccd1 vccd1 o_data1[14] sky130_fd_sc_hd__buf_2
X_9237_ clknet_leaf_20_i_clk _0381_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6449_ reg_data\[2\]\[1\] _1021_ _1064_ _1105_ reg_data\[11\]\[1\] vssd1 vssd1 vccd1
+ vccd1 _3010_ sky130_fd_sc_hd__a32o_1
X_9168_ clknet_leaf_22_i_clk _0312_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_8119_ _3869_ reg_data\[13\]\[5\] _3963_ vssd1 vssd1 vccd1 vccd1 _3969_ sky130_fd_sc_hd__mux2_1
X_9099_ clknet_leaf_27_i_clk _0243_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_2_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5820_ _1115_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__buf_2
X_5751_ _1021_ vssd1 vssd1 vccd1 vccd1 _2336_ sky130_fd_sc_hd__clkbuf_4
X_8470_ _4143_ vssd1 vssd1 vccd1 vccd1 _4155_ sky130_fd_sc_hd__buf_4
X_4702_ reg_data\[0\]\[4\] _1070_ _1318_ _1319_ _1320_ vssd1 vssd1 vccd1 vccd1 _1321_
+ sky130_fd_sc_hd__a2111o_1
X_5682_ reg_data\[0\]\[20\] _1775_ _2266_ _2267_ _2268_ vssd1 vssd1 vccd1 vccd1 _2269_
+ sky130_fd_sc_hd__a2111o_1
X_7421_ _3581_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__clkbuf_1
X_4633_ _1056_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__buf_4
X_4564_ _1171_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__buf_2
X_7352_ reg_data\[3\]\[14\] _3158_ _3540_ vssd1 vssd1 vccd1 vccd1 _3545_ sky130_fd_sc_hd__mux2_1
X_6303_ reg_data\[6\]\[30\] _2555_ _1270_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__and3_1
X_7283_ _3508_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__clkbuf_1
X_6234_ reg_data\[27\]\[29\] _2392_ _2800_ _2801_ _2802_ vssd1 vssd1 vccd1 vccd1 _2803_
+ sky130_fd_sc_hd__a2111o_1
X_4495_ _1021_ _1117_ _1094_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__and3_4
X_9022_ clknet_leaf_74_i_clk _0166_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6165_ reg_data\[30\]\[28\] _2524_ _1919_ vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__and3_1
X_6096_ reg_data\[23\]\[26\] _2440_ _2441_ reg_data\[19\]\[26\] vssd1 vssd1 vccd1
+ vccd1 _2670_ sky130_fd_sc_hd__a22o_1
X_5116_ reg_data\[0\]\[11\] _1070_ _1717_ _1719_ _1720_ vssd1 vssd1 vccd1 vccd1 _1721_
+ sky130_fd_sc_hd__a2111o_1
X_5047_ reg_data\[21\]\[10\] _1480_ _1240_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__and3_1
X_9855_ clknet_leaf_24_i_clk rs2_mux\[2\] vssd1 vssd1 vccd1 vccd1 rs2\[2\] sky130_fd_sc_hd__dfxtp_1
X_9786_ clknet_leaf_55_i_clk rdata1\[2\] vssd1 vssd1 vccd1 vccd1 r_data1\[2\] sky130_fd_sc_hd__dfxtp_1
X_8806_ reg_data\[11\]\[8\] i_data[8] _4324_ vssd1 vssd1 vccd1 vccd1 _4333_ sky130_fd_sc_hd__mux2_1
X_6998_ _3355_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__clkbuf_1
X_5949_ reg_data\[6\]\[24\] _2207_ _2323_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__and3_1
X_8737_ _4296_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__clkbuf_1
X_8668_ reg_data\[19\]\[7\] _3143_ _4252_ vssd1 vssd1 vccd1 vccd1 _4260_ sky130_fd_sc_hd__mux2_1
X_7619_ _3676_ vssd1 vssd1 vccd1 vccd1 _3688_ sky130_fd_sc_hd__buf_4
X_8599_ _4223_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__clkbuf_1
X_7970_ i_data[10] vssd1 vssd1 vccd1 vccd1 _3879_ sky130_fd_sc_hd__buf_2
X_6921_ _3212_ reg_data\[10\]\[5\] _3309_ vssd1 vssd1 vccd1 vccd1 _3315_ sky130_fd_sc_hd__mux2_1
X_6852_ _3277_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__clkbuf_1
X_9640_ clknet_leaf_49_i_clk _0784_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_5803_ _1080_ vssd1 vssd1 vccd1 vccd1 _2386_ sky130_fd_sc_hd__clkbuf_4
X_9571_ clknet_leaf_60_i_clk _0715_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8522_ reg_data\[1\]\[2\] _3133_ _4180_ vssd1 vssd1 vccd1 vccd1 _4183_ sky130_fd_sc_hd__mux2_1
X_6783_ _3231_ reg_data\[22\]\[14\] _3223_ vssd1 vssd1 vccd1 vccd1 _3232_ sky130_fd_sc_hd__mux2_1
X_5734_ reg_data\[18\]\[21\] _2261_ _2090_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__and3_1
X_8453_ _4146_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__clkbuf_1
X_5665_ reg_data\[26\]\[19\] _1849_ _1850_ reg_data\[29\]\[19\] vssd1 vssd1 vccd1
+ vccd1 _2253_ sky130_fd_sc_hd__a22o_1
X_8384_ _3861_ reg_data\[17\]\[1\] _4108_ vssd1 vssd1 vccd1 vccd1 _4110_ sky130_fd_sc_hd__mux2_1
X_7404_ _3572_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__clkbuf_1
X_4616_ reg_data\[22\]\[3\] _1039_ _1236_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__and3_1
X_5596_ reg_data\[12\]\[18\] _1960_ _2016_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__and3_1
X_7335_ reg_data\[3\]\[6\] _3141_ _3529_ vssd1 vssd1 vccd1 vccd1 _3536_ sky130_fd_sc_hd__mux2_1
X_4547_ reg_data\[18\]\[2\] _1166_ _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__and3_1
X_4478_ _1100_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__buf_4
X_7266_ _3499_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
X_6217_ reg_data\[25\]\[29\] _2370_ _2783_ _2784_ _2785_ vssd1 vssd1 vccd1 vccd1 _2786_
+ sky130_fd_sc_hd__a2111o_1
X_9005_ clknet_leaf_27_i_clk _0149_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_7197_ _3462_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__clkbuf_1
X_6148_ reg_data\[7\]\[27\] _2433_ _2717_ _2718_ _2719_ vssd1 vssd1 vccd1 vccd1 _2720_
+ sky130_fd_sc_hd__a2111o_1
X_6079_ reg_data\[22\]\[26\] _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__and3_1
X_9907_ clknet_leaf_57_i_clk _0977_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_9838_ clknet_leaf_39_i_clk rdata2\[22\] vssd1 vssd1 vccd1 vccd1 r_data2\[22\] sky130_fd_sc_hd__dfxtp_1
X_9769_ clknet_leaf_57_i_clk _0913_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_20_i_clk clknet_3_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_35_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5450_ reg_data\[7\]\[16\] _1780_ _2042_ _2043_ _2044_ vssd1 vssd1 vccd1 vccd1 _2045_
+ sky130_fd_sc_hd__a2111o_1
X_4401_ _1026_ vssd1 vssd1 vccd1 vccd1 rs1_mux\[1\] sky130_fd_sc_hd__inv_2
X_5381_ reg_data\[30\]\[15\] _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__and3_1
X_7120_ reg_data\[7\]\[1\] _3131_ _3420_ vssd1 vssd1 vccd1 vccd1 _3422_ sky130_fd_sc_hd__mux2_1
X_7051_ _3204_ reg_data\[8\]\[1\] _3383_ vssd1 vssd1 vccd1 vccd1 _3385_ sky130_fd_sc_hd__mux2_1
X_6002_ reg_data\[18\]\[25\] _2261_ _2090_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__and3_1
X_7953_ _3867_ reg_data\[9\]\[4\] _3859_ vssd1 vssd1 vccd1 vccd1 _3868_ sky130_fd_sc_hd__mux2_1
X_6904_ _3304_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__clkbuf_1
X_7884_ _3214_ reg_data\[28\]\[6\] _3822_ vssd1 vssd1 vccd1 vccd1 _3829_ sky130_fd_sc_hd__mux2_1
X_6835_ _3266_ reg_data\[22\]\[31\] _3201_ vssd1 vssd1 vccd1 vccd1 _3267_ sky130_fd_sc_hd__mux2_1
X_9623_ clknet_leaf_43_i_clk _0767_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_9554_ clknet_leaf_17_i_clk _0698_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6766_ i_data[9] vssd1 vssd1 vccd1 vccd1 _3220_ sky130_fd_sc_hd__buf_2
X_8505_ _4173_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__clkbuf_1
X_5717_ reg_data\[12\]\[20\] _1960_ _2016_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__and3_1
X_9485_ clknet_leaf_29_i_clk _0629_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6697_ reg_data\[4\]\[20\] _3170_ _3171_ vssd1 vssd1 vccd1 vccd1 _3172_ sky130_fd_sc_hd__mux2_1
X_8436_ _3913_ reg_data\[17\]\[26\] _4130_ vssd1 vssd1 vccd1 vccd1 _4137_ sky130_fd_sc_hd__mux2_1
X_5648_ reg_data\[3\]\[19\] _1815_ _2232_ _2233_ _2235_ vssd1 vssd1 vccd1 vccd1 _2236_
+ sky130_fd_sc_hd__a2111o_1
X_8367_ _4100_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__clkbuf_1
X_5579_ _2161_ _2165_ _2167_ _2169_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__or4_1
X_8298_ _4063_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__clkbuf_1
X_7318_ _3526_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__clkbuf_1
X_7249_ _3489_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkbuf_1
X_4950_ reg_data\[24\]\[8\] _1127_ _1130_ reg_data\[28\]\[8\] _1560_ vssd1 vssd1 vccd1
+ vccd1 _1561_ sky130_fd_sc_hd__a221o_1
X_4881_ reg_data\[14\]\[7\] _1381_ _1090_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__and3_1
X_6620_ _3116_ vssd1 vssd1 vccd1 vccd1 o_data2[30] sky130_fd_sc_hd__buf_2
X_6551_ _3079_ vssd1 vssd1 vccd1 vccd1 o_data1[30] sky130_fd_sc_hd__buf_2
X_5502_ reg_data\[6\]\[17\] _1600_ _1716_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__and3_1
X_9270_ clknet_leaf_39_i_clk _0414_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6482_ reg_data\[24\]\[1\] _1224_ _1227_ reg_data\[28\]\[1\] _3041_ vssd1 vssd1 vccd1
+ vccd1 _3042_ sky130_fd_sc_hd__a221o_1
X_8221_ _3903_ reg_data\[14\]\[21\] _4021_ vssd1 vssd1 vccd1 vccd1 _4023_ sky130_fd_sc_hd__mux2_1
X_5433_ _2028_ vssd1 vssd1 vccd1 vccd1 rdata2\[15\] sky130_fd_sc_hd__clkbuf_1
X_8152_ _3986_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__clkbuf_1
X_5364_ reg_data\[7\]\[14\] _1827_ _1957_ _1959_ _1961_ vssd1 vssd1 vccd1 vccd1 _1962_
+ sky130_fd_sc_hd__a2111o_1
X_7103_ _3256_ reg_data\[8\]\[26\] _3405_ vssd1 vssd1 vccd1 vccd1 _3412_ sky130_fd_sc_hd__mux2_1
X_8083_ _3949_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__clkbuf_1
X_5295_ reg_data\[13\]\[13\] _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__and3_1
X_7034_ _3374_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__clkbuf_1
X_8985_ clknet_leaf_12_i_clk _0129_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_7936_ _3266_ reg_data\[28\]\[31\] _3821_ vssd1 vssd1 vccd1 vccd1 _3856_ sky130_fd_sc_hd__mux2_1
X_7867_ _3266_ reg_data\[27\]\[31\] _3784_ vssd1 vssd1 vccd1 vccd1 _3819_ sky130_fd_sc_hd__mux2_1
X_6818_ _3255_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__clkbuf_1
X_9606_ clknet_leaf_51_i_clk _0750_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_7798_ _3782_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__clkbuf_1
X_6749_ _3208_ reg_data\[22\]\[3\] _3202_ vssd1 vssd1 vccd1 vccd1 _3209_ sky130_fd_sc_hd__mux2_1
X_9537_ clknet_leaf_5_i_clk _0681_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_9468_ clknet_leaf_10_i_clk _0612_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_8419_ _3896_ reg_data\[17\]\[18\] _4119_ vssd1 vssd1 vccd1 vccd1 _4128_ sky130_fd_sc_hd__mux2_1
X_9399_ clknet_leaf_43_i_clk _0543_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5080_ reg_data\[20\]\[10\] _1629_ _1180_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__and3_1
X_8770_ _3907_ reg_data\[29\]\[23\] _4310_ vssd1 vssd1 vccd1 vccd1 _4314_ sky130_fd_sc_hd__mux2_1
X_5982_ reg_data\[13\]\[24\] _2183_ _2299_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__and3_1
X_7721_ _3256_ reg_data\[25\]\[26\] _3735_ vssd1 vssd1 vccd1 vccd1 _3742_ sky130_fd_sc_hd__mux2_1
X_4933_ reg_data\[3\]\[8\] _1054_ _1541_ _1542_ _1543_ vssd1 vssd1 vccd1 vccd1 _1544_
+ sky130_fd_sc_hd__a2111o_1
X_7652_ _3705_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__clkbuf_1
X_4864_ _1477_ vssd1 vssd1 vccd1 vccd1 rdata2\[6\] sky130_fd_sc_hd__clkbuf_1
X_7583_ _3668_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__clkbuf_1
X_6603_ r_data2\[22\] _3105_ vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__and2_1
X_4795_ reg_data\[13\]\[5\] _1186_ _1191_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__and3_1
X_9322_ clknet_leaf_40_i_clk _0466_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6534_ r_data1\[22\] _3068_ vssd1 vssd1 vccd1 vccd1 _3071_ sky130_fd_sc_hd__and2_1
X_6465_ reg_data\[3\]\[1\] _1157_ _3022_ _3023_ _3024_ vssd1 vssd1 vccd1 vccd1 _3025_
+ sky130_fd_sc_hd__a2111o_1
X_9253_ clknet_leaf_57_i_clk _0397_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5416_ reg_data\[5\]\[15\] _1824_ _1954_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__and3_1
X_8204_ _3886_ reg_data\[14\]\[13\] _4010_ vssd1 vssd1 vccd1 vccd1 _4014_ sky130_fd_sc_hd__mux2_1
X_6396_ reg_data\[1\]\[0\] _1103_ _1108_ _1110_ reg_data\[15\]\[0\] vssd1 vssd1 vccd1
+ vccd1 _2959_ sky130_fd_sc_hd__a32o_1
X_9184_ clknet_leaf_2_i_clk _0328_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_5347_ reg_data\[17\]\[14\] _1509_ _1275_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__and3_1
X_8135_ _3977_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__clkbuf_1
X_5278_ reg_data\[26\]\[13\] _1805_ _1806_ reg_data\[29\]\[13\] vssd1 vssd1 vccd1
+ vccd1 _1879_ sky130_fd_sc_hd__a22o_1
X_8066_ _3940_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__clkbuf_1
X_7017_ _3365_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__clkbuf_1
X_8968_ clknet_leaf_54_i_clk _0112_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_7919_ _3847_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__clkbuf_1
X_8899_ clknet_leaf_64_i_clk _0043_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_4580_ _1000_ _1147_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__and2_2
X_6250_ reg_data\[4\]\[29\] _1175_ _1342_ vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__and3_1
X_6181_ reg_data\[16\]\[28\] _2405_ _2406_ reg_data\[9\]\[28\] vssd1 vssd1 vccd1 vccd1
+ _2752_ sky130_fd_sc_hd__a22o_1
X_5201_ _1129_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__clkbuf_4
X_5132_ _1736_ vssd1 vssd1 vccd1 vccd1 rdata1\[11\] sky130_fd_sc_hd__clkbuf_1
X_5063_ reg_data\[23\]\[10\] _1099_ _1101_ reg_data\[19\]\[10\] vssd1 vssd1 vccd1
+ vccd1 _1670_ sky130_fd_sc_hd__a22o_1
X_9871_ clknet_leaf_58_i_clk _0941_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8822_ _4341_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__clkbuf_1
X_5965_ reg_data\[26\]\[24\] _2411_ _2412_ reg_data\[29\]\[24\] vssd1 vssd1 vccd1
+ vccd1 _2544_ sky130_fd_sc_hd__a22o_1
X_8753_ _3890_ reg_data\[29\]\[15\] _4299_ vssd1 vssd1 vccd1 vccd1 _4305_ sky130_fd_sc_hd__mux2_1
X_5896_ reg_data\[7\]\[23\] _2386_ _2474_ _2475_ _2476_ vssd1 vssd1 vccd1 vccd1 _2477_
+ sky130_fd_sc_hd__a2111o_1
X_7704_ _3239_ reg_data\[25\]\[18\] _3724_ vssd1 vssd1 vccd1 vccd1 _3733_ sky130_fd_sc_hd__mux2_1
X_8684_ _4268_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__clkbuf_1
X_4916_ reg_data\[2\]\[7\] _1002_ _1295_ _1296_ reg_data\[11\]\[7\] vssd1 vssd1 vccd1
+ vccd1 _1528_ sky130_fd_sc_hd__a32o_1
X_7635_ _3696_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__clkbuf_1
X_4847_ reg_data\[4\]\[6\] _1460_ _1407_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__and3_1
X_9305_ clknet_leaf_9_i_clk _0449_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_4778_ _1394_ vssd1 vssd1 vccd1 vccd1 rdata1\[5\] sky130_fd_sc_hd__dlymetal6s2s_1
X_7566_ _3659_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__clkbuf_1
X_7497_ _3622_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__clkbuf_1
X_6517_ r_data1\[14\] _3057_ vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__and2_1
X_9236_ clknet_leaf_21_i_clk _0380_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6448_ reg_data\[23\]\[1\] _1098_ _1100_ reg_data\[19\]\[1\] vssd1 vssd1 vccd1 vccd1
+ _3009_ sky130_fd_sc_hd__a22o_1
X_9167_ clknet_leaf_30_i_clk _0311_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6379_ reg_data\[21\]\[0\] _1058_ _1044_ vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__and3_1
X_8118_ _3968_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__clkbuf_1
X_9098_ clknet_leaf_42_i_clk _0242_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8049_ _3931_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__clkbuf_1
X_5750_ reg_data\[2\]\[21\] _2219_ _1790_ _1791_ reg_data\[11\]\[21\] vssd1 vssd1
+ vccd1 vccd1 _2335_ sky130_fd_sc_hd__a32o_1
X_5681_ reg_data\[5\]\[20\] _2097_ _1925_ vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__and3_1
X_4701_ reg_data\[5\]\[4\] _1076_ _1250_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__and3_1
X_4632_ _1071_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__clkbuf_4
X_7420_ _3231_ reg_data\[20\]\[14\] _3576_ vssd1 vssd1 vccd1 vccd1 _3581_ sky130_fd_sc_hd__mux2_1
X_4563_ _1184_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__clkbuf_4
X_7351_ _3544_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__clkbuf_1
X_6302_ reg_data\[3\]\[30\] _2421_ _2865_ _2866_ _2867_ vssd1 vssd1 vccd1 vccd1 _2868_
+ sky130_fd_sc_hd__a2111o_1
X_4494_ rs1_mux\[0\] _1026_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__nor2_1
X_7282_ reg_data\[5\]\[13\] _3156_ _3504_ vssd1 vssd1 vccd1 vccd1 _3508_ sky130_fd_sc_hd__mux2_1
X_6233_ reg_data\[1\]\[29\] _2336_ _2399_ _2400_ reg_data\[15\]\[29\] vssd1 vssd1
+ vccd1 vccd1 _2802_ sky130_fd_sc_hd__a32o_1
X_9021_ clknet_leaf_70_i_clk _0165_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6164_ reg_data\[18\]\[28\] _2261_ _1063_ vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__and3_1
X_6095_ _2656_ _2660_ _2664_ _2668_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__or4_2
X_5115_ reg_data\[5\]\[11\] _1490_ _1250_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__and3_1
X_5046_ reg_data\[17\]\[10\] _1042_ _1238_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__and3_1
X_9854_ clknet_leaf_24_i_clk rs2_mux\[1\] vssd1 vssd1 vccd1 vccd1 rs2\[1\] sky130_fd_sc_hd__dfxtp_1
X_9785_ clknet_leaf_56_i_clk rdata1\[1\] vssd1 vssd1 vccd1 vccd1 r_data1\[1\] sky130_fd_sc_hd__dfxtp_1
X_8805_ _4332_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__clkbuf_1
X_6997_ reg_data\[0\]\[9\] _3147_ _3345_ vssd1 vssd1 vccd1 vccd1 _3355_ sky130_fd_sc_hd__mux2_1
X_5948_ reg_data\[3\]\[24\] _2376_ _2523_ _2525_ _2526_ vssd1 vssd1 vccd1 vccd1 _2527_
+ sky130_fd_sc_hd__a2111o_1
X_8736_ _3873_ reg_data\[29\]\[7\] _4288_ vssd1 vssd1 vccd1 vccd1 _4296_ sky130_fd_sc_hd__mux2_1
X_5879_ reg_data\[22\]\[23\] _2143_ _2256_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__and3_1
X_8667_ _4259_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__clkbuf_1
X_7618_ _3687_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__clkbuf_1
X_8598_ _3871_ reg_data\[12\]\[6\] _4216_ vssd1 vssd1 vccd1 vccd1 _4223_ sky130_fd_sc_hd__mux2_1
X_7549_ _3650_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__clkbuf_1
X_9219_ clknet_leaf_64_i_clk _0363_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6920_ _3314_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__clkbuf_1
X_6851_ reg_data\[2\]\[5\] _3139_ _3271_ vssd1 vssd1 vccd1 vccd1 _3277_ sky130_fd_sc_hd__mux2_1
X_5802_ reg_data\[0\]\[22\] _2381_ _2382_ _2383_ _2384_ vssd1 vssd1 vccd1 vccd1 _2385_
+ sky130_fd_sc_hd__a2111o_1
X_9570_ clknet_leaf_60_i_clk _0714_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6782_ i_data[14] vssd1 vssd1 vccd1 vccd1 _3231_ sky130_fd_sc_hd__buf_2
X_8521_ _4182_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__clkbuf_1
X_5733_ reg_data\[25\]\[21\] _1764_ _2315_ _2316_ _2317_ vssd1 vssd1 vccd1 vccd1 _2318_
+ sky130_fd_sc_hd__a2111o_1
X_8452_ _3861_ reg_data\[18\]\[1\] _4144_ vssd1 vssd1 vccd1 vccd1 _4146_ sky130_fd_sc_hd__mux2_1
X_5664_ reg_data\[8\]\[19\] _1841_ _1842_ reg_data\[10\]\[19\] _2251_ vssd1 vssd1
+ vccd1 vccd1 _2252_ sky130_fd_sc_hd__a221o_1
X_4615_ _1047_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__buf_2
X_8383_ _4109_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__clkbuf_1
X_5595_ reg_data\[14\]\[18\] _1693_ _1958_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__and3_1
X_7403_ _3214_ reg_data\[20\]\[6\] _3565_ vssd1 vssd1 vccd1 vccd1 _3572_ sky130_fd_sc_hd__mux2_1
X_7334_ _3535_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__clkbuf_1
X_4546_ _1167_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__buf_4
X_4477_ _1097_ _1051_ _1052_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__and3_4
X_7265_ reg_data\[5\]\[5\] _3139_ _3493_ vssd1 vssd1 vccd1 vccd1 _3499_ sky130_fd_sc_hd__mux2_1
X_6216_ reg_data\[21\]\[29\] _1058_ _2087_ vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__and3_1
X_9004_ clknet_leaf_27_i_clk _0148_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_7196_ reg_data\[6\]\[5\] _3139_ _3456_ vssd1 vssd1 vccd1 vccd1 _3462_ sky130_fd_sc_hd__mux2_1
X_6147_ reg_data\[13\]\[27\] _2562_ _1191_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__and3_1
X_6078_ _2652_ vssd1 vssd1 vccd1 vccd1 rdata1\[26\] sky130_fd_sc_hd__clkbuf_1
X_9906_ clknet_leaf_56_i_clk _0976_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_5029_ reg_data\[13\]\[9\] _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__and3_1
X_9837_ clknet_leaf_39_i_clk rdata2\[21\] vssd1 vssd1 vccd1 vccd1 r_data2\[21\] sky130_fd_sc_hd__dfxtp_1
X_9768_ clknet_leaf_56_i_clk _0912_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_1_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_8719_ _4286_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__clkbuf_1
X_9699_ clknet_leaf_60_i_clk _0843_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_4400_ _1025_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__buf_2
X_5380_ reg_data\[18\]\[15\] _1656_ _1483_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__and3_1
X_7050_ _3384_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__clkbuf_1
X_6001_ reg_data\[25\]\[25\] _2370_ _2575_ _2576_ _2577_ vssd1 vssd1 vccd1 vccd1 _2578_
+ sky130_fd_sc_hd__a2111o_1
X_7952_ i_data[4] vssd1 vssd1 vccd1 vccd1 _3867_ sky130_fd_sc_hd__clkbuf_4
X_6903_ reg_data\[2\]\[30\] _3191_ _3270_ vssd1 vssd1 vccd1 vccd1 _3304_ sky130_fd_sc_hd__mux2_1
X_9622_ clknet_leaf_43_i_clk _0766_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_7883_ _3828_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__clkbuf_1
X_6834_ i_data[31] vssd1 vssd1 vccd1 vccd1 _3266_ sky130_fd_sc_hd__clkbuf_4
X_9553_ clknet_leaf_17_i_clk _0697_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6765_ _3219_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__clkbuf_1
X_8504_ _3913_ reg_data\[18\]\[26\] _4166_ vssd1 vssd1 vccd1 vccd1 _4173_ sky130_fd_sc_hd__mux2_1
X_9484_ clknet_leaf_29_i_clk _0628_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5716_ reg_data\[14\]\[20\] _2301_ _1958_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__and3_1
X_8435_ _4136_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__clkbuf_1
X_6696_ _3128_ vssd1 vssd1 vccd1 vccd1 _3171_ sky130_fd_sc_hd__buf_4
X_5647_ reg_data\[20\]\[19\] _2234_ _1743_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__and3_1
X_8366_ _3911_ reg_data\[16\]\[25\] _4094_ vssd1 vssd1 vccd1 vccd1 _4100_ sky130_fd_sc_hd__mux2_1
X_5578_ reg_data\[24\]\[18\] _1803_ _1804_ reg_data\[28\]\[18\] _2168_ vssd1 vssd1
+ vccd1 vccd1 _2169_ sky130_fd_sc_hd__a221o_1
X_8297_ _3911_ reg_data\[15\]\[25\] _4057_ vssd1 vssd1 vccd1 vccd1 _4063_ sky130_fd_sc_hd__mux2_1
X_4529_ _1005_ _1013_ rs2_mux\[2\] _0993_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__and4b_2
X_7317_ reg_data\[5\]\[30\] _3191_ _3492_ vssd1 vssd1 vccd1 vccd1 _3526_ sky130_fd_sc_hd__mux2_1
X_7248_ reg_data\[6\]\[30\] _3191_ _3455_ vssd1 vssd1 vccd1 vccd1 _3489_ sky130_fd_sc_hd__mux2_1
X_7179_ _3452_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__clkbuf_1
X_4880_ reg_data\[13\]\[7\] _1253_ _1087_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__and3_1
X_6550_ r_data1\[30\] _3045_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__and2_1
X_5501_ reg_data\[3\]\[17\] _1770_ _2091_ _2092_ _2093_ vssd1 vssd1 vccd1 vccd1 _2094_
+ sky130_fd_sc_hd__a2111o_1
X_6481_ reg_data\[26\]\[1\] _1229_ _1231_ reg_data\[29\]\[1\] vssd1 vssd1 vccd1 vccd1
+ _3041_ sky130_fd_sc_hd__a22o_1
X_8220_ _4022_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__clkbuf_1
X_5432_ _2019_ _2023_ _2025_ _2027_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__or4_1
X_8151_ _3900_ reg_data\[13\]\[20\] _3985_ vssd1 vssd1 vccd1 vccd1 _3986_ sky130_fd_sc_hd__mux2_1
X_5363_ reg_data\[12\]\[14\] _1960_ _1226_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__and3_1
X_7102_ _3411_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__clkbuf_1
X_8082_ _3900_ reg_data\[30\]\[20\] _3948_ vssd1 vssd1 vccd1 vccd1 _3949_ sky130_fd_sc_hd__mux2_1
X_5294_ reg_data\[0\]\[13\] _1821_ _1891_ _1892_ _1893_ vssd1 vssd1 vccd1 vccd1 _1894_
+ sky130_fd_sc_hd__a2111o_1
X_7033_ reg_data\[0\]\[26\] _3183_ _3367_ vssd1 vssd1 vccd1 vccd1 _3374_ sky130_fd_sc_hd__mux2_1
X_8984_ clknet_leaf_13_i_clk _0128_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_7935_ _3855_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__clkbuf_1
X_7866_ _3818_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__clkbuf_1
X_6817_ _3254_ reg_data\[22\]\[25\] _3244_ vssd1 vssd1 vccd1 vccd1 _3255_ sky130_fd_sc_hd__mux2_1
X_9605_ clknet_leaf_52_i_clk _0749_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_7797_ _3264_ reg_data\[26\]\[30\] _3748_ vssd1 vssd1 vccd1 vccd1 _3782_ sky130_fd_sc_hd__mux2_1
X_9536_ clknet_leaf_5_i_clk _0680_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6748_ i_data[3] vssd1 vssd1 vccd1 vccd1 _3208_ sky130_fd_sc_hd__buf_2
X_6679_ _3159_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__clkbuf_1
X_9467_ clknet_leaf_4_i_clk _0611_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_9398_ clknet_leaf_39_i_clk _0542_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_8418_ _4127_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__clkbuf_1
X_8349_ _3894_ reg_data\[16\]\[17\] _4083_ vssd1 vssd1 vccd1 vccd1 _4091_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_34_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_49_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_3_4__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5981_ reg_data\[0\]\[24\] _2427_ _2556_ _2557_ _2558_ vssd1 vssd1 vccd1 vccd1 _2559_
+ sky130_fd_sc_hd__a2111o_1
X_7720_ _3741_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__clkbuf_1
X_4932_ reg_data\[20\]\[8\] _1062_ _1315_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__and3_1
X_7651_ _3254_ reg_data\[24\]\[25\] _3699_ vssd1 vssd1 vccd1 vccd1 _3705_ sky130_fd_sc_hd__mux2_1
X_6602_ _3107_ vssd1 vssd1 vccd1 vccd1 o_data2[21] sky130_fd_sc_hd__buf_2
X_4863_ _1468_ _1472_ _1474_ _1476_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__or4_1
X_7582_ reg_data\[23\]\[25\] _3181_ _3662_ vssd1 vssd1 vccd1 vccd1 _3668_ sky130_fd_sc_hd__mux2_1
X_4794_ reg_data\[0\]\[5\] _1174_ _1406_ _1408_ _1409_ vssd1 vssd1 vccd1 vccd1 _1410_
+ sky130_fd_sc_hd__a2111o_1
X_6533_ _3070_ vssd1 vssd1 vccd1 vccd1 o_data1[21] sky130_fd_sc_hd__buf_2
X_9321_ clknet_leaf_41_i_clk _0465_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6464_ reg_data\[20\]\[1\] _1150_ _1283_ vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__and3_1
X_9252_ clknet_leaf_60_i_clk _0396_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8203_ _4013_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__clkbuf_1
X_5415_ reg_data\[4\]\[15\] _1460_ _1407_ vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__and3_1
X_6395_ reg_data\[2\]\[0\] _1021_ _1064_ _1105_ reg_data\[11\]\[0\] vssd1 vssd1 vccd1
+ vccd1 _2958_ sky130_fd_sc_hd__a32o_1
X_9183_ clknet_leaf_1_i_clk _0327_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8134_ _3884_ reg_data\[13\]\[12\] _3974_ vssd1 vssd1 vccd1 vccd1 _3977_ sky130_fd_sc_hd__mux2_1
X_5346_ reg_data\[21\]\[14\] _1883_ _1943_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__and3_1
X_5277_ reg_data\[8\]\[13\] _1797_ _1798_ reg_data\[10\]\[13\] _1877_ vssd1 vssd1
+ vccd1 vccd1 _1878_ sky130_fd_sc_hd__a221o_1
X_8065_ _3884_ reg_data\[30\]\[12\] _3937_ vssd1 vssd1 vccd1 vccd1 _3940_ sky130_fd_sc_hd__mux2_1
X_7016_ reg_data\[0\]\[18\] _3166_ _3356_ vssd1 vssd1 vccd1 vccd1 _3365_ sky130_fd_sc_hd__mux2_1
X_8967_ clknet_leaf_51_i_clk _0111_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_7918_ _3248_ reg_data\[28\]\[22\] _3844_ vssd1 vssd1 vccd1 vccd1 _3847_ sky130_fd_sc_hd__mux2_1
X_8898_ clknet_leaf_63_i_clk _0042_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_7849_ _3248_ reg_data\[27\]\[22\] _3807_ vssd1 vssd1 vccd1 vccd1 _3810_ sky130_fd_sc_hd__mux2_1
X_9519_ clknet_leaf_23_i_clk _0663_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6180_ reg_data\[27\]\[28\] _2392_ _2748_ _2749_ _2750_ vssd1 vssd1 vccd1 vccd1 _2751_
+ sky130_fd_sc_hd__a2111o_1
X_5200_ _1126_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__clkbuf_4
X_5131_ _1726_ _1731_ _1733_ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__or4_1
X_5062_ _1655_ _1660_ _1664_ _1668_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__or4_1
X_9870_ clknet_leaf_62_i_clk _0940_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8821_ reg_data\[11\]\[15\] i_data[15] _4335_ vssd1 vssd1 vccd1 vccd1 _4341_ sky130_fd_sc_hd__mux2_1
X_8752_ _4304_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__clkbuf_1
X_5964_ reg_data\[8\]\[24\] _2403_ _2404_ reg_data\[10\]\[24\] _2542_ vssd1 vssd1
+ vccd1 vccd1 _2543_ sky130_fd_sc_hd__a221o_1
X_7703_ _3732_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__clkbuf_1
X_5895_ reg_data\[12\]\[23\] _2214_ _1128_ vssd1 vssd1 vccd1 vccd1 _2476_ sky130_fd_sc_hd__and3_1
X_4915_ reg_data\[23\]\[7\] _1206_ _1209_ reg_data\[19\]\[7\] vssd1 vssd1 vccd1 vccd1
+ _1527_ sky130_fd_sc_hd__a22o_1
X_8683_ reg_data\[19\]\[14\] _3158_ _4263_ vssd1 vssd1 vccd1 vccd1 _4268_ sky130_fd_sc_hd__mux2_1
X_7634_ _3237_ reg_data\[24\]\[17\] _3688_ vssd1 vssd1 vccd1 vccd1 _3696_ sky130_fd_sc_hd__mux2_1
X_4846_ _0999_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__clkbuf_4
X_7565_ reg_data\[23\]\[17\] _3164_ _3651_ vssd1 vssd1 vccd1 vccd1 _3659_ sky130_fd_sc_hd__mux2_1
X_9304_ clknet_leaf_9_i_clk _0448_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_4777_ _1385_ _1389_ _1391_ _1393_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__or4_1
X_6516_ _3061_ vssd1 vssd1 vccd1 vccd1 o_data1[13] sky130_fd_sc_hd__buf_2
X_7496_ _3237_ reg_data\[21\]\[17\] _3614_ vssd1 vssd1 vccd1 vccd1 _3622_ sky130_fd_sc_hd__mux2_1
X_9235_ clknet_leaf_21_i_clk _0379_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6447_ _2995_ _2999_ _3003_ _3007_ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__or4_2
X_9166_ clknet_leaf_29_i_clk _0310_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6378_ reg_data\[17\]\[0\] _1055_ _1040_ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__and3_1
X_5329_ reg_data\[14\]\[14\] _1867_ _1379_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__and3_1
X_8117_ _3867_ reg_data\[13\]\[4\] _3963_ vssd1 vssd1 vccd1 vccd1 _3968_ sky130_fd_sc_hd__mux2_1
X_9097_ clknet_leaf_42_i_clk _0241_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_8048_ _3867_ reg_data\[30\]\[4\] _3926_ vssd1 vssd1 vccd1 vccd1 _3931_ sky130_fd_sc_hd__mux2_1
X_5680_ reg_data\[4\]\[20\] _1718_ _1863_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__and3_1
X_4700_ reg_data\[4\]\[4\] _1074_ _1248_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__and3_1
X_4631_ reg_data\[0\]\[3\] _1070_ _1247_ _1249_ _1251_ vssd1 vssd1 vccd1 vccd1 _1252_
+ sky130_fd_sc_hd__a2111o_1
X_4562_ _1171_ _1183_ _1156_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__and3_2
X_7350_ reg_data\[3\]\[13\] _3156_ _3540_ vssd1 vssd1 vccd1 vccd1 _3544_ sky130_fd_sc_hd__mux2_1
X_6301_ reg_data\[20\]\[30\] _1150_ _1283_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__and3_1
X_4493_ _1115_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__clkbuf_4
X_7281_ _3507_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__clkbuf_1
X_6232_ reg_data\[2\]\[29\] _1021_ _2396_ _2397_ reg_data\[11\]\[29\] vssd1 vssd1
+ vccd1 vccd1 _2801_ sky130_fd_sc_hd__a32o_1
X_9020_ clknet_leaf_74_i_clk _0164_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6163_ reg_data\[25\]\[28\] _2370_ _2731_ _2732_ _2733_ vssd1 vssd1 vccd1 vccd1 _2734_
+ sky130_fd_sc_hd__a2111o_1
X_6094_ reg_data\[7\]\[26\] _2433_ _2665_ _2666_ _2667_ vssd1 vssd1 vccd1 vccd1 _2668_
+ sky130_fd_sc_hd__a2111o_1
X_5114_ reg_data\[4\]\[11\] _1718_ _1248_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__and3_1
X_5045_ reg_data\[22\]\[10\] _1536_ _1651_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__and3_1
X_9853_ clknet_leaf_24_i_clk rs2_mux\[0\] vssd1 vssd1 vccd1 vccd1 rs2\[0\] sky130_fd_sc_hd__dfxtp_1
X_9784_ clknet_leaf_56_i_clk rdata1\[0\] vssd1 vssd1 vccd1 vccd1 r_data1\[0\] sky130_fd_sc_hd__dfxtp_1
X_8804_ reg_data\[11\]\[7\] i_data[7] _4324_ vssd1 vssd1 vccd1 vccd1 _4332_ sky130_fd_sc_hd__mux2_1
X_6996_ _3354_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__clkbuf_1
X_5947_ reg_data\[30\]\[24\] _2204_ _1254_ vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__and3_1
X_8735_ _4295_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__clkbuf_1
X_8666_ reg_data\[19\]\[6\] _3141_ _4252_ vssd1 vssd1 vccd1 vccd1 _4259_ sky130_fd_sc_hd__mux2_1
X_5878_ _2459_ vssd1 vssd1 vccd1 vccd1 rdata2\[22\] sky130_fd_sc_hd__clkbuf_1
X_7617_ _3220_ reg_data\[24\]\[9\] _3677_ vssd1 vssd1 vccd1 vccd1 _3687_ sky130_fd_sc_hd__mux2_1
X_4829_ reg_data\[1\]\[6\] _1022_ _1109_ _1111_ reg_data\[15\]\[6\] vssd1 vssd1 vccd1
+ vccd1 _1444_ sky130_fd_sc_hd__a32o_1
X_8597_ _4222_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__clkbuf_1
X_7548_ reg_data\[23\]\[9\] _3147_ _3640_ vssd1 vssd1 vccd1 vccd1 _3650_ sky130_fd_sc_hd__mux2_1
X_7479_ _3220_ reg_data\[21\]\[9\] _3603_ vssd1 vssd1 vccd1 vccd1 _3613_ sky130_fd_sc_hd__mux2_1
X_9218_ clknet_leaf_66_i_clk _0362_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_9149_ clknet_leaf_3_i_clk _0293_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6850_ _3276_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkbuf_1
X_5801_ reg_data\[5\]\[22\] _2097_ _1925_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__and3_1
X_6781_ _3230_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__clkbuf_1
X_5732_ reg_data\[21\]\[21\] _2086_ _2087_ vssd1 vssd1 vccd1 vccd1 _2317_ sky130_fd_sc_hd__and3_1
X_8520_ reg_data\[1\]\[1\] _3131_ _4180_ vssd1 vssd1 vccd1 vccd1 _4182_ sky130_fd_sc_hd__mux2_1
X_8451_ _4145_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__clkbuf_1
X_5663_ reg_data\[16\]\[19\] _1843_ _1844_ reg_data\[9\]\[19\] vssd1 vssd1 vccd1 vccd1
+ _2251_ sky130_fd_sc_hd__a22o_1
X_8382_ _3857_ reg_data\[17\]\[0\] _4108_ vssd1 vssd1 vccd1 vccd1 _4109_ sky130_fd_sc_hd__mux2_1
X_5594_ reg_data\[13\]\[18\] _2183_ _1576_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__and3_1
X_4614_ _1235_ vssd1 vssd1 vccd1 vccd1 rdata2\[2\] sky130_fd_sc_hd__dlymetal6s2s_1
X_7402_ _3571_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__clkbuf_1
X_4545_ rs2_mux\[0\] _1006_ _1010_ _1013_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__and4bb_4
X_7333_ reg_data\[3\]\[5\] _3139_ _3529_ vssd1 vssd1 vccd1 vccd1 _3535_ sky130_fd_sc_hd__mux2_1
X_9003_ clknet_leaf_43_i_clk _0147_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_4476_ _1098_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__buf_4
X_7264_ _3498_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
X_6215_ reg_data\[17\]\[29\] _2372_ _1040_ vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__and3_1
X_7195_ _3461_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__clkbuf_1
X_6146_ reg_data\[12\]\[27\] _2301_ _1187_ vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__and3_1
X_6077_ _2643_ _2647_ _2649_ _2651_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__or4_1
X_9905_ clknet_leaf_56_i_clk _0975_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_5028_ reg_data\[0\]\[9\] _1174_ _1633_ _1634_ _1635_ vssd1 vssd1 vccd1 vccd1 _1636_
+ sky130_fd_sc_hd__a2111o_1
X_9836_ clknet_leaf_40_i_clk rdata2\[20\] vssd1 vssd1 vccd1 vccd1 r_data2\[20\] sky130_fd_sc_hd__dfxtp_1
X_6979_ reg_data\[0\]\[0\] _3118_ _3345_ vssd1 vssd1 vccd1 vccd1 _3346_ sky130_fd_sc_hd__mux2_1
X_9767_ clknet_leaf_56_i_clk _0911_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8718_ reg_data\[19\]\[31\] _3193_ _4251_ vssd1 vssd1 vccd1 vccd1 _4286_ sky130_fd_sc_hd__mux2_1
X_9698_ clknet_leaf_60_i_clk _0842_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8649_ _4249_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__clkbuf_1
X_6000_ reg_data\[21\]\[25\] _2086_ _2087_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__and3_1
X_7951_ _3866_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__clkbuf_1
X_6902_ _3303_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__clkbuf_1
X_7882_ _3212_ reg_data\[28\]\[5\] _3822_ vssd1 vssd1 vccd1 vccd1 _3828_ sky130_fd_sc_hd__mux2_1
X_9621_ clknet_leaf_32_i_clk _0765_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6833_ _3265_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__clkbuf_1
X_9552_ clknet_leaf_19_i_clk _0696_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6764_ _3218_ reg_data\[22\]\[8\] _3202_ vssd1 vssd1 vccd1 vccd1 _3219_ sky130_fd_sc_hd__mux2_1
X_8503_ _4172_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__clkbuf_1
X_5715_ _1171_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__clkbuf_4
X_9483_ clknet_leaf_27_i_clk _0627_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6695_ i_data[20] vssd1 vssd1 vccd1 vccd1 _3170_ sky130_fd_sc_hd__clkbuf_4
X_8434_ _3911_ reg_data\[17\]\[25\] _4130_ vssd1 vssd1 vccd1 vccd1 _4136_ sky130_fd_sc_hd__mux2_1
X_5646_ _1138_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__clkbuf_4
X_8365_ _4099_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__clkbuf_1
X_5577_ reg_data\[26\]\[18\] _1805_ _1806_ reg_data\[29\]\[18\] vssd1 vssd1 vccd1
+ vccd1 _2168_ sky130_fd_sc_hd__a22o_1
X_8296_ _4062_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__clkbuf_1
X_7316_ _3525_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__clkbuf_1
X_4528_ _1138_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__buf_2
X_7247_ _3488_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__clkbuf_1
X_4459_ _1071_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__buf_2
X_7178_ reg_data\[7\]\[29\] _3189_ _3442_ vssd1 vssd1 vccd1 vccd1 _3452_ sky130_fd_sc_hd__mux2_1
X_6129_ reg_data\[26\]\[27\] _2411_ _2412_ reg_data\[29\]\[27\] vssd1 vssd1 vccd1
+ vccd1 _2702_ sky130_fd_sc_hd__a22o_1
X_9819_ clknet_leaf_60_i_clk rdata2\[3\] vssd1 vssd1 vccd1 vccd1 r_data2\[3\] sky130_fd_sc_hd__dfxtp_1
X_5500_ reg_data\[20\]\[17\] _1597_ _2035_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__and3_1
X_6480_ reg_data\[8\]\[1\] _1213_ _1216_ reg_data\[10\]\[1\] _3039_ vssd1 vssd1 vccd1
+ vccd1 _3040_ sky130_fd_sc_hd__a221o_1
X_5431_ reg_data\[24\]\[15\] _1847_ _1848_ reg_data\[28\]\[15\] _2026_ vssd1 vssd1
+ vccd1 vccd1 _2027_ sky130_fd_sc_hd__a221o_1
X_8150_ _3962_ vssd1 vssd1 vccd1 vccd1 _3985_ sky130_fd_sc_hd__buf_4
X_5362_ _1000_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__buf_2
X_7101_ _3254_ reg_data\[8\]\[25\] _3405_ vssd1 vssd1 vccd1 vccd1 _3411_ sky130_fd_sc_hd__mux2_1
X_8081_ _3925_ vssd1 vssd1 vccd1 vccd1 _3948_ sky130_fd_sc_hd__buf_4
X_7032_ _3373_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_0_i_clk clknet_3_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5293_ reg_data\[5\]\[13\] _1824_ _1285_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__and3_1
X_8983_ clknet_leaf_43_i_clk _0127_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_7934_ _3264_ reg_data\[28\]\[30\] _3821_ vssd1 vssd1 vccd1 vccd1 _3855_ sky130_fd_sc_hd__mux2_1
X_7865_ _3264_ reg_data\[27\]\[30\] _3784_ vssd1 vssd1 vccd1 vccd1 _3818_ sky130_fd_sc_hd__mux2_1
X_7796_ _3781_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__clkbuf_1
X_6816_ i_data[25] vssd1 vssd1 vccd1 vccd1 _3254_ sky130_fd_sc_hd__clkbuf_4
X_9604_ clknet_leaf_62_i_clk _0748_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_9535_ clknet_leaf_4_i_clk _0679_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6747_ _3207_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__clkbuf_1
X_9466_ clknet_leaf_10_i_clk _0610_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6678_ reg_data\[4\]\[14\] _3158_ _3150_ vssd1 vssd1 vccd1 vccd1 _3159_ sky130_fd_sc_hd__mux2_1
X_9397_ clknet_leaf_37_i_clk _0541_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_8417_ _3894_ reg_data\[17\]\[17\] _4119_ vssd1 vssd1 vccd1 vccd1 _4127_ sky130_fd_sc_hd__mux2_1
X_5629_ reg_data\[23\]\[19\] _1787_ _1788_ reg_data\[19\]\[19\] vssd1 vssd1 vccd1
+ vccd1 _2218_ sky130_fd_sc_hd__a22o_1
X_8348_ _4090_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__clkbuf_1
X_8279_ _4053_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__clkbuf_1
X_5980_ reg_data\[5\]\[24\] _2430_ _1338_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__and3_1
X_4931_ reg_data\[30\]\[8\] _1312_ _1313_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__and3_1
X_7650_ _3704_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__clkbuf_1
X_4862_ reg_data\[24\]\[6\] _1225_ _1228_ reg_data\[28\]\[6\] _1475_ vssd1 vssd1 vccd1
+ vccd1 _1476_ sky130_fd_sc_hd__a221o_1
X_6601_ r_data2\[21\] _3105_ vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__and2_1
X_7581_ _3667_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__clkbuf_1
X_4793_ reg_data\[5\]\[5\] _1179_ _1285_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__and3_1
X_9320_ clknet_leaf_49_i_clk _0464_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6532_ r_data1\[21\] _3068_ vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__and2_1
X_6463_ reg_data\[30\]\[1\] _1146_ _1163_ vssd1 vssd1 vccd1 vccd1 _3023_ sky130_fd_sc_hd__and3_1
X_9251_ clknet_leaf_60_i_clk _0395_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_9182_ clknet_leaf_2_i_clk _0326_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8202_ _3884_ reg_data\[14\]\[12\] _4010_ vssd1 vssd1 vccd1 vccd1 _4013_ sky130_fd_sc_hd__mux2_1
X_5414_ reg_data\[6\]\[15\] _1951_ _1632_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__and3_1
X_6394_ reg_data\[23\]\[0\] _1098_ _1100_ reg_data\[19\]\[0\] vssd1 vssd1 vccd1 vccd1
+ _2957_ sky130_fd_sc_hd__a22o_1
X_8133_ _3976_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__clkbuf_1
X_5345_ _1144_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__buf_4
X_5276_ reg_data\[16\]\[13\] _1799_ _1800_ reg_data\[9\]\[13\] vssd1 vssd1 vccd1 vccd1
+ _1877_ sky130_fd_sc_hd__a22o_1
X_8064_ _3939_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__clkbuf_1
X_7015_ _3364_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__clkbuf_1
X_8966_ clknet_leaf_50_i_clk _0110_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_7917_ _3846_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__clkbuf_1
X_8897_ clknet_leaf_66_i_clk _0041_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_7848_ _3809_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__clkbuf_1
X_7779_ _3246_ reg_data\[26\]\[21\] _3771_ vssd1 vssd1 vccd1 vccd1 _3773_ sky130_fd_sc_hd__mux2_1
X_9518_ clknet_leaf_23_i_clk _0662_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_9449_ clknet_leaf_62_i_clk _0593_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_5130_ reg_data\[24\]\[11\] _1127_ _1130_ reg_data\[28\]\[11\] _1734_ vssd1 vssd1
+ vccd1 vccd1 _1735_ sky130_fd_sc_hd__a221o_1
X_5061_ reg_data\[7\]\[10\] _1081_ _1665_ _1666_ _1667_ vssd1 vssd1 vccd1 vccd1 _1668_
+ sky130_fd_sc_hd__a2111o_1
X_8820_ _4340_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__clkbuf_1
X_5963_ reg_data\[16\]\[24\] _2405_ _2406_ reg_data\[9\]\[24\] vssd1 vssd1 vccd1 vccd1
+ _2542_ sky130_fd_sc_hd__a22o_1
X_8751_ _3888_ reg_data\[29\]\[14\] _4299_ vssd1 vssd1 vccd1 vccd1 _4304_ sky130_fd_sc_hd__mux2_1
X_4914_ _1512_ _1517_ _1521_ _1525_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__or4_1
X_7702_ _3237_ reg_data\[25\]\[17\] _3724_ vssd1 vssd1 vccd1 vccd1 _3732_ sky130_fd_sc_hd__mux2_1
X_5894_ reg_data\[14\]\[23\] _1986_ _1090_ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__and3_1
X_8682_ _4267_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__clkbuf_1
X_7633_ _3695_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__clkbuf_1
X_4845_ reg_data\[6\]\[6\] _1347_ _1152_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__and3_1
X_4776_ reg_data\[24\]\[5\] _1127_ _1130_ reg_data\[28\]\[5\] _1392_ vssd1 vssd1 vccd1
+ vccd1 _1393_ sky130_fd_sc_hd__a221o_1
X_7564_ _3658_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__clkbuf_1
X_9303_ clknet_leaf_43_i_clk _0447_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6515_ r_data1\[13\] _3057_ vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_33_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_7495_ _3621_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__clkbuf_1
X_9234_ clknet_leaf_30_i_clk _0378_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6446_ reg_data\[7\]\[1\] _1080_ _3004_ _3005_ _3006_ vssd1 vssd1 vccd1 vccd1 _3007_
+ sky130_fd_sc_hd__a2111o_1
X_9165_ clknet_leaf_29_i_clk _0309_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6377_ reg_data\[22\]\[0\] _1097_ _1047_ vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__and3_1
X_5328_ reg_data\[0\]\[14\] _1775_ _1923_ _1924_ _1926_ vssd1 vssd1 vccd1 vccd1 _1927_
+ sky130_fd_sc_hd__a2111o_1
X_9096_ clknet_leaf_48_i_clk _0240_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_8116_ _3967_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_48_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_8047_ _3930_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__clkbuf_1
X_5259_ reg_data\[20\]\[13\] _1597_ _1315_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__and3_1
X_8949_ clknet_leaf_36_i_clk _0093_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_4630_ reg_data\[5\]\[3\] _1076_ _1250_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__and3_1
X_6300_ reg_data\[30\]\[30\] _1146_ _1163_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__and3_1
X_4561_ _1010_ rs2_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__nor2_1
X_4492_ _1089_ _1094_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__and3_4
X_7280_ reg_data\[5\]\[12\] _3154_ _3504_ vssd1 vssd1 vccd1 vccd1 _3507_ sky130_fd_sc_hd__mux2_1
X_6231_ reg_data\[23\]\[29\] _2393_ _2394_ reg_data\[19\]\[29\] vssd1 vssd1 vccd1
+ vccd1 _2800_ sky130_fd_sc_hd__a22o_1
X_6162_ reg_data\[21\]\[28\] _1058_ _2087_ vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__and3_1
X_5113_ _1071_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__clkbuf_4
X_6093_ reg_data\[12\]\[26\] _2562_ _1289_ vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__and3_1
X_9921_ clknet_leaf_43_i_clk _0991_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5044_ _1047_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__clkbuf_4
X_9852_ clknet_leaf_20_i_clk rs1_mux\[4\] vssd1 vssd1 vccd1 vccd1 rs1\[4\] sky130_fd_sc_hd__dfxtp_1
X_8803_ _4331_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__clkbuf_1
X_9783_ clknet_leaf_39_i_clk _0927_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6995_ reg_data\[0\]\[8\] _3145_ _3345_ vssd1 vssd1 vccd1 vccd1 _3354_ sky130_fd_sc_hd__mux2_1
X_5946_ reg_data\[20\]\[24\] _2524_ _1060_ vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__and3_1
X_8734_ _3871_ reg_data\[29\]\[6\] _4288_ vssd1 vssd1 vccd1 vccd1 _4295_ sky130_fd_sc_hd__mux2_1
X_5877_ _2438_ _2446_ _2452_ _2458_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__or4_1
X_8665_ _4258_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__clkbuf_1
X_4828_ reg_data\[2\]\[6\] _1103_ _1104_ _1106_ reg_data\[11\]\[6\] vssd1 vssd1 vccd1
+ vccd1 _1443_ sky130_fd_sc_hd__a32o_1
X_7616_ _3686_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__clkbuf_1
X_8596_ _3869_ reg_data\[12\]\[5\] _4216_ vssd1 vssd1 vccd1 vccd1 _4222_ sky130_fd_sc_hd__mux2_1
X_7547_ _3649_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__clkbuf_1
X_4759_ reg_data\[4\]\[5\] _1074_ _1248_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__and3_1
X_7478_ _3612_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__clkbuf_1
X_6429_ _2982_ _2986_ _2988_ _2990_ vssd1 vssd1 vccd1 vccd1 _2991_ sky130_fd_sc_hd__or4_2
X_9217_ clknet_leaf_6_i_clk _0361_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_9148_ clknet_leaf_11_i_clk _0292_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_9079_ clknet_leaf_14_i_clk _0223_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5800_ reg_data\[4\]\[22\] _2325_ _1863_ vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__and3_1
X_6780_ _3229_ reg_data\[22\]\[13\] _3223_ vssd1 vssd1 vccd1 vccd1 _3230_ sky130_fd_sc_hd__mux2_1
X_5731_ reg_data\[17\]\[21\] _1766_ _1708_ vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__and3_1
X_8450_ _3857_ reg_data\[18\]\[0\] _4144_ vssd1 vssd1 vccd1 vccd1 _4145_ sky130_fd_sc_hd__mux2_1
X_5662_ reg_data\[27\]\[19\] _1833_ _2247_ _2248_ _2249_ vssd1 vssd1 vccd1 vccd1 _2250_
+ sky130_fd_sc_hd__a2111o_1
X_5593_ _1171_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__clkbuf_4
X_8381_ _4107_ vssd1 vssd1 vccd1 vccd1 _4108_ sky130_fd_sc_hd__buf_4
X_4613_ _1196_ _1211_ _1223_ _1234_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__or4_1
X_7401_ _3212_ reg_data\[20\]\[5\] _3565_ vssd1 vssd1 vccd1 vccd1 _3571_ sky130_fd_sc_hd__mux2_1
X_4544_ _1138_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__buf_2
X_7332_ _3534_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__clkbuf_1
X_7263_ reg_data\[5\]\[4\] _3137_ _3493_ vssd1 vssd1 vccd1 vccd1 _3498_ sky130_fd_sc_hd__mux2_1
X_6214_ reg_data\[22\]\[29\] _1097_ _2256_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__and3_1
X_4475_ _1097_ _1079_ _1052_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__and3_4
X_9002_ clknet_leaf_42_i_clk _0146_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_7194_ reg_data\[6\]\[4\] _3137_ _3456_ vssd1 vssd1 vccd1 vccd1 _3461_ sky130_fd_sc_hd__mux2_1
X_6145_ reg_data\[14\]\[27\] _2183_ _1164_ vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__and3_1
X_6076_ reg_data\[24\]\[26\] _2409_ _2410_ reg_data\[28\]\[26\] _2650_ vssd1 vssd1
+ vccd1 vccd1 _2651_ sky130_fd_sc_hd__a221o_1
X_9904_ clknet_leaf_57_i_clk _0974_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_5027_ reg_data\[5\]\[9\] _1179_ _1285_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__and3_1
X_9835_ clknet_leaf_52_i_clk rdata2\[19\] vssd1 vssd1 vccd1 vccd1 r_data2\[19\] sky130_fd_sc_hd__dfxtp_1
X_9766_ clknet_leaf_55_i_clk _0910_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6978_ _3344_ vssd1 vssd1 vccd1 vccd1 _3345_ sky130_fd_sc_hd__buf_4
X_8717_ _4285_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__clkbuf_1
X_5929_ reg_data\[2\]\[23\] _2443_ _2507_ _2508_ reg_data\[11\]\[23\] vssd1 vssd1
+ vccd1 vccd1 _2509_ sky130_fd_sc_hd__a32o_1
X_9697_ clknet_leaf_1_i_clk _0841_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_8648_ _3921_ reg_data\[12\]\[30\] _4215_ vssd1 vssd1 vccd1 vccd1 _4249_ sky130_fd_sc_hd__mux2_1
X_8579_ _4212_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__clkbuf_1
X_7950_ _3865_ reg_data\[9\]\[3\] _3859_ vssd1 vssd1 vccd1 vccd1 _3866_ sky130_fd_sc_hd__mux2_1
X_6901_ reg_data\[2\]\[29\] _3189_ _3293_ vssd1 vssd1 vccd1 vccd1 _3303_ sky130_fd_sc_hd__mux2_1
X_7881_ _3827_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__clkbuf_1
X_9620_ clknet_leaf_32_i_clk _0764_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6832_ _3264_ reg_data\[22\]\[30\] _3201_ vssd1 vssd1 vccd1 vccd1 _3265_ sky130_fd_sc_hd__mux2_1
X_9551_ clknet_leaf_22_i_clk _0695_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6763_ i_data[8] vssd1 vssd1 vccd1 vccd1 _3218_ sky130_fd_sc_hd__clkbuf_4
X_8502_ _3911_ reg_data\[18\]\[25\] _4166_ vssd1 vssd1 vccd1 vccd1 _4172_ sky130_fd_sc_hd__mux2_1
X_5714_ reg_data\[13\]\[20\] _2183_ _2299_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__and3_1
X_6694_ _3169_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__clkbuf_1
X_9482_ clknet_leaf_44_i_clk _0626_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8433_ _4135_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__clkbuf_1
X_5645_ reg_data\[30\]\[19\] _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__and3_1
X_8364_ _3909_ reg_data\[16\]\[24\] _4094_ vssd1 vssd1 vccd1 vccd1 _4099_ sky130_fd_sc_hd__mux2_1
X_5576_ reg_data\[8\]\[18\] _1797_ _1798_ reg_data\[10\]\[18\] _2166_ vssd1 vssd1
+ vccd1 vccd1 _2167_ sky130_fd_sc_hd__a221o_1
X_8295_ _3909_ reg_data\[15\]\[24\] _4057_ vssd1 vssd1 vccd1 vccd1 _4062_ sky130_fd_sc_hd__mux2_1
X_7315_ reg_data\[5\]\[29\] _3189_ _3515_ vssd1 vssd1 vccd1 vccd1 _3525_ sky130_fd_sc_hd__mux2_1
X_4527_ reg_data\[17\]\[2\] _1146_ _1148_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__and3_1
X_7246_ reg_data\[6\]\[29\] _3189_ _3478_ vssd1 vssd1 vccd1 vccd1 _3488_ sky130_fd_sc_hd__mux2_1
X_4458_ _1080_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__clkbuf_4
X_7177_ _3451_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__clkbuf_1
X_6128_ reg_data\[8\]\[27\] _2403_ _2404_ reg_data\[10\]\[27\] _2700_ vssd1 vssd1
+ vccd1 vccd1 _2701_ sky130_fd_sc_hd__a221o_1
X_4389_ i_rs1[0] i_rs1[2] i_rs1[3] i_rs1[1] vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__or4_1
X_6059_ reg_data\[3\]\[26\] _2376_ _2631_ _2632_ _2633_ vssd1 vssd1 vccd1 vccd1 _2634_
+ sky130_fd_sc_hd__a2111o_1
X_9818_ clknet_leaf_54_i_clk rdata2\[2\] vssd1 vssd1 vccd1 vccd1 r_data2\[2\] sky130_fd_sc_hd__dfxtp_1
X_9749_ clknet_leaf_16_i_clk _0893_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_5430_ reg_data\[26\]\[15\] _1849_ _1850_ reg_data\[29\]\[15\] vssd1 vssd1 vccd1
+ vccd1 _2026_ sky130_fd_sc_hd__a22o_1
X_5361_ reg_data\[14\]\[14\] _1693_ _1958_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__and3_1
X_7100_ _3410_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__clkbuf_1
X_8080_ _3947_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__clkbuf_1
X_5292_ reg_data\[4\]\[13\] _1460_ _1407_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__and3_1
X_7031_ reg_data\[0\]\[25\] _3181_ _3367_ vssd1 vssd1 vccd1 vccd1 _3373_ sky130_fd_sc_hd__mux2_1
X_8982_ clknet_leaf_43_i_clk _0126_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_7933_ _3854_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__clkbuf_1
X_7864_ _3817_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__clkbuf_1
X_7795_ _3262_ reg_data\[26\]\[29\] _3771_ vssd1 vssd1 vccd1 vccd1 _3781_ sky130_fd_sc_hd__mux2_1
X_6815_ _3253_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__clkbuf_1
X_9603_ clknet_leaf_62_i_clk _0747_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_9534_ clknet_leaf_4_i_clk _0678_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6746_ _3206_ reg_data\[22\]\[2\] _3202_ vssd1 vssd1 vccd1 vccd1 _3207_ sky130_fd_sc_hd__mux2_1
X_9465_ clknet_leaf_11_i_clk _0609_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6677_ i_data[14] vssd1 vssd1 vccd1 vccd1 _3158_ sky130_fd_sc_hd__clkbuf_4
X_9396_ clknet_leaf_32_i_clk _0540_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_5628_ _2201_ _2206_ _2211_ _2216_ vssd1 vssd1 vccd1 vccd1 _2217_ sky130_fd_sc_hd__or4_2
X_8416_ _4126_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__clkbuf_1
X_5559_ reg_data\[20\]\[18\] _1597_ _2035_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__and3_1
X_8347_ _3892_ reg_data\[16\]\[16\] _4083_ vssd1 vssd1 vccd1 vccd1 _4090_ sky130_fd_sc_hd__mux2_1
X_8278_ _3892_ reg_data\[15\]\[16\] _4046_ vssd1 vssd1 vccd1 vccd1 _4053_ sky130_fd_sc_hd__mux2_1
X_7229_ _3479_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__clkbuf_1
X_4930_ reg_data\[18\]\[8\] _1055_ _1483_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__and3_1
X_4861_ reg_data\[26\]\[6\] _1230_ _1232_ reg_data\[29\]\[6\] vssd1 vssd1 vccd1 vccd1
+ _1475_ sky130_fd_sc_hd__a22o_1
X_6600_ _3106_ vssd1 vssd1 vccd1 vccd1 o_data2[20] sky130_fd_sc_hd__buf_2
X_7580_ reg_data\[23\]\[24\] _3179_ _3662_ vssd1 vssd1 vccd1 vccd1 _3667_ sky130_fd_sc_hd__mux2_1
X_4792_ reg_data\[4\]\[5\] _1177_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__and3_1
X_6531_ _3069_ vssd1 vssd1 vccd1 vccd1 o_data1[20] sky130_fd_sc_hd__buf_2
X_6462_ reg_data\[18\]\[1\] _1143_ _1167_ vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__and3_1
X_9250_ clknet_leaf_60_i_clk _0394_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6393_ _2943_ _2947_ _2951_ _2955_ vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__or4_2
X_9181_ clknet_leaf_1_i_clk _0325_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_5413_ reg_data\[3\]\[15\] _1815_ _2004_ _2007_ _2008_ vssd1 vssd1 vccd1 vccd1 _2009_
+ sky130_fd_sc_hd__a2111o_1
X_8201_ _4012_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__clkbuf_1
X_5344_ reg_data\[22\]\[14\] _1679_ _1622_ vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__and3_1
X_8132_ _3882_ reg_data\[13\]\[11\] _3974_ vssd1 vssd1 vccd1 vccd1 _3976_ sky130_fd_sc_hd__mux2_1
X_5275_ reg_data\[27\]\[13\] _1786_ _1873_ _1874_ _1875_ vssd1 vssd1 vccd1 vccd1 _1876_
+ sky130_fd_sc_hd__a2111o_1
X_8063_ _3882_ reg_data\[30\]\[11\] _3937_ vssd1 vssd1 vccd1 vccd1 _3939_ sky130_fd_sc_hd__mux2_1
X_7014_ reg_data\[0\]\[17\] _3164_ _3356_ vssd1 vssd1 vccd1 vccd1 _3364_ sky130_fd_sc_hd__mux2_1
X_8965_ clknet_leaf_51_i_clk _0109_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8896_ clknet_leaf_67_i_clk _0040_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7916_ _3246_ reg_data\[28\]\[21\] _3844_ vssd1 vssd1 vccd1 vccd1 _3846_ sky130_fd_sc_hd__mux2_1
X_7847_ _3246_ reg_data\[27\]\[21\] _3807_ vssd1 vssd1 vccd1 vccd1 _3809_ sky130_fd_sc_hd__mux2_1
X_7778_ _3772_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__clkbuf_1
X_9517_ clknet_leaf_25_i_clk _0661_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6729_ i_data[31] vssd1 vssd1 vccd1 vccd1 _3193_ sky130_fd_sc_hd__buf_4
X_9448_ clknet_leaf_51_i_clk _0592_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_9379_ clknet_leaf_60_i_clk _0523_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_5060_ reg_data\[13\]\[10\] _1608_ _1257_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__and3_1
X_5962_ reg_data\[27\]\[24\] _2392_ _2538_ _2539_ _2540_ vssd1 vssd1 vccd1 vccd1 _2541_
+ sky130_fd_sc_hd__a2111o_1
X_8750_ _4303_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__clkbuf_1
X_4913_ reg_data\[7\]\[7\] _1185_ _1522_ _1523_ _1524_ vssd1 vssd1 vccd1 vccd1 _1525_
+ sky130_fd_sc_hd__a2111o_1
X_7701_ _3731_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__clkbuf_1
X_5893_ reg_data\[13\]\[23\] _2473_ _1087_ vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__and3_1
X_8681_ reg_data\[19\]\[13\] _3156_ _4263_ vssd1 vssd1 vccd1 vccd1 _4267_ sky130_fd_sc_hd__mux2_1
X_7632_ _3235_ reg_data\[24\]\[16\] _3688_ vssd1 vssd1 vccd1 vccd1 _3695_ sky130_fd_sc_hd__mux2_1
X_4844_ reg_data\[3\]\[6\] _1158_ _1455_ _1456_ _1457_ vssd1 vssd1 vccd1 vccd1 _1458_
+ sky130_fd_sc_hd__a2111o_1
X_4775_ reg_data\[26\]\[5\] _1132_ _1134_ reg_data\[29\]\[5\] vssd1 vssd1 vccd1 vccd1
+ _1392_ sky130_fd_sc_hd__a22o_1
X_7563_ reg_data\[23\]\[16\] _3162_ _3651_ vssd1 vssd1 vccd1 vccd1 _3658_ sky130_fd_sc_hd__mux2_1
X_9302_ clknet_leaf_38_i_clk _0446_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6514_ _3060_ vssd1 vssd1 vccd1 vccd1 o_data1[12] sky130_fd_sc_hd__buf_2
X_9233_ clknet_leaf_22_i_clk _0377_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_7494_ _3235_ reg_data\[21\]\[16\] _3614_ vssd1 vssd1 vccd1 vccd1 _3621_ sky130_fd_sc_hd__mux2_1
X_6445_ reg_data\[13\]\[1\] _1076_ _1087_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__and3_1
X_6376_ _2939_ vssd1 vssd1 vccd1 vccd1 rdata2\[31\] sky130_fd_sc_hd__clkbuf_1
X_9164_ clknet_leaf_27_i_clk _0308_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5327_ reg_data\[5\]\[14\] _1490_ _1925_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__and3_1
X_9095_ clknet_leaf_48_i_clk _0239_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8115_ _3865_ reg_data\[13\]\[3\] _3963_ vssd1 vssd1 vccd1 vccd1 _3967_ sky130_fd_sc_hd__mux2_1
X_8046_ _3865_ reg_data\[30\]\[3\] _3926_ vssd1 vssd1 vccd1 vccd1 _3930_ sky130_fd_sc_hd__mux2_1
X_5258_ reg_data\[30\]\[13\] _1312_ _1313_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__and3_1
X_5189_ reg_data\[2\]\[12\] _1613_ _1790_ _1791_ reg_data\[11\]\[12\] vssd1 vssd1
+ vccd1 vccd1 _1792_ sky130_fd_sc_hd__a32o_1
X_8948_ clknet_leaf_37_i_clk _0092_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_8879_ clknet_leaf_29_i_clk _0023_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_4560_ reg_data\[0\]\[2\] _1174_ _1176_ _1178_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_
+ sky130_fd_sc_hd__a2111o_1
X_4491_ rs1_mux\[0\] rs1_mux\[1\] vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__nor2_1
X_6230_ _2786_ _2790_ _2794_ _2798_ vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__or4_4
X_6161_ reg_data\[17\]\[28\] _2372_ _1040_ vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__and3_1
X_5112_ reg_data\[6\]\[11\] _1600_ _1716_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__and3_1
X_6092_ reg_data\[14\]\[26\] _2301_ _1344_ vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__and3_1
X_9920_ clknet_leaf_43_i_clk _0990_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_5043_ _1650_ vssd1 vssd1 vccd1 vccd1 rdata2\[9\] sky130_fd_sc_hd__clkbuf_1
X_9851_ clknet_leaf_24_i_clk rs1_mux\[3\] vssd1 vssd1 vccd1 vccd1 rs1\[3\] sky130_fd_sc_hd__dfxtp_1
X_8802_ reg_data\[11\]\[6\] i_data[6] _4324_ vssd1 vssd1 vccd1 vccd1 _4331_ sky130_fd_sc_hd__mux2_1
X_9782_ clknet_leaf_39_i_clk _0926_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6994_ _3353_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__clkbuf_1
X_5945_ _1038_ vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__buf_2
X_8733_ _4294_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__clkbuf_1
X_5876_ reg_data\[24\]\[22\] _2453_ _2454_ reg_data\[28\]\[22\] _2457_ vssd1 vssd1
+ vccd1 vccd1 _2458_ sky130_fd_sc_hd__a221o_1
X_8664_ reg_data\[19\]\[5\] _3139_ _4252_ vssd1 vssd1 vccd1 vccd1 _4258_ sky130_fd_sc_hd__mux2_1
X_4827_ reg_data\[23\]\[6\] _1099_ _1101_ reg_data\[19\]\[6\] vssd1 vssd1 vccd1 vccd1
+ _1442_ sky130_fd_sc_hd__a22o_1
X_7615_ _3218_ reg_data\[24\]\[8\] _3677_ vssd1 vssd1 vccd1 vccd1 _3686_ sky130_fd_sc_hd__mux2_1
X_8595_ _4221_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__clkbuf_1
X_7546_ reg_data\[23\]\[8\] _3145_ _3640_ vssd1 vssd1 vccd1 vccd1 _3649_ sky130_fd_sc_hd__mux2_1
X_4758_ reg_data\[6\]\[5\] _1072_ _1048_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__and3_1
X_7477_ _3218_ reg_data\[21\]\[8\] _3603_ vssd1 vssd1 vccd1 vccd1 _3612_ sky130_fd_sc_hd__mux2_1
X_4689_ reg_data\[21\]\[4\] _1042_ _1044_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__and3_1
X_6428_ reg_data\[24\]\[0\] _1224_ _1227_ reg_data\[28\]\[0\] _2989_ vssd1 vssd1 vccd1
+ vccd1 _2990_ sky130_fd_sc_hd__a221o_1
X_9216_ clknet_leaf_66_i_clk _0360_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_9147_ clknet_leaf_4_i_clk _0291_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6359_ reg_data\[4\]\[31\] _1175_ _1342_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__and3_1
X_9078_ clknet_leaf_16_i_clk _0222_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_8029_ i_data[29] vssd1 vssd1 vccd1 vccd1 _3919_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_32_i_clk clknet_3_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5730_ reg_data\[22\]\[21\] _2143_ _2256_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__and3_1
X_5661_ reg_data\[1\]\[19\] _1904_ _1905_ reg_data\[15\]\[19\] vssd1 vssd1 vccd1 vccd1
+ _2249_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_47_i_clk clknet_3_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_7400_ _3570_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__clkbuf_1
X_5592_ reg_data\[0\]\[18\] _1821_ _2179_ _2180_ _2181_ vssd1 vssd1 vccd1 vccd1 _2182_
+ sky130_fd_sc_hd__a2111o_1
X_8380_ _3601_ _4070_ vssd1 vssd1 vccd1 vccd1 _4107_ sky130_fd_sc_hd__nand2_2
X_4612_ reg_data\[24\]\[2\] _1225_ _1228_ reg_data\[28\]\[2\] _1233_ vssd1 vssd1 vccd1
+ vccd1 _1234_ sky130_fd_sc_hd__a221o_1
X_4543_ reg_data\[30\]\[2\] _1162_ _1164_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__and3_1
X_7331_ reg_data\[3\]\[4\] _3137_ _3529_ vssd1 vssd1 vccd1 vccd1 _3534_ sky130_fd_sc_hd__mux2_1
X_7262_ _3497_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__clkbuf_1
X_6213_ _2782_ vssd1 vssd1 vccd1 vccd1 rdata2\[28\] sky130_fd_sc_hd__clkbuf_1
X_4474_ _1017_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__buf_2
X_9001_ clknet_leaf_42_i_clk _0145_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_7193_ _3460_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__clkbuf_1
X_6144_ reg_data\[0\]\[27\] _2427_ _2713_ _2714_ _2715_ vssd1 vssd1 vccd1 vccd1 _2716_
+ sky130_fd_sc_hd__a2111o_1
X_6075_ reg_data\[26\]\[26\] _2411_ _2412_ reg_data\[29\]\[26\] vssd1 vssd1 vccd1
+ vccd1 _2650_ sky130_fd_sc_hd__a22o_1
X_9903_ clknet_leaf_59_i_clk _0973_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5026_ reg_data\[4\]\[9\] _1460_ _1407_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__and3_1
X_9834_ clknet_leaf_50_i_clk rdata2\[18\] vssd1 vssd1 vccd1 vccd1 r_data2\[18\] sky130_fd_sc_hd__dfxtp_1
X_6977_ _3127_ _3269_ vssd1 vssd1 vccd1 vccd1 _3344_ sky130_fd_sc_hd__nor2_4
X_9765_ clknet_leaf_57_i_clk _0909_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8716_ reg_data\[19\]\[30\] _3191_ _4251_ vssd1 vssd1 vccd1 vccd1 _4285_ sky130_fd_sc_hd__mux2_1
X_5928_ _1200_ vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__buf_4
X_9696_ clknet_leaf_75_i_clk _0840_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8647_ _4248_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__clkbuf_1
X_5859_ _1208_ vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__buf_2
X_8578_ reg_data\[1\]\[29\] _3189_ _4202_ vssd1 vssd1 vccd1 vccd1 _4212_ sky130_fd_sc_hd__mux2_1
X_7529_ _3639_ vssd1 vssd1 vccd1 vccd1 _3640_ sky130_fd_sc_hd__buf_4
X_6900_ _3302_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__clkbuf_1
X_7880_ _3210_ reg_data\[28\]\[4\] _3822_ vssd1 vssd1 vccd1 vccd1 _3827_ sky130_fd_sc_hd__mux2_1
X_6831_ i_data[30] vssd1 vssd1 vccd1 vccd1 _3264_ sky130_fd_sc_hd__clkbuf_4
X_9550_ clknet_leaf_23_i_clk _0694_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_8501_ _4171_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__clkbuf_1
X_6762_ _3217_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__clkbuf_1
X_5713_ _1190_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__clkbuf_4
X_6693_ reg_data\[4\]\[19\] _3168_ _3150_ vssd1 vssd1 vccd1 vccd1 _3169_ sky130_fd_sc_hd__mux2_1
X_9481_ clknet_leaf_44_i_clk _0625_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_8432_ _3909_ reg_data\[17\]\[24\] _4130_ vssd1 vssd1 vccd1 vccd1 _4135_ sky130_fd_sc_hd__mux2_1
X_5644_ reg_data\[18\]\[19\] _1816_ _2120_ vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__and3_1
X_8363_ _4098_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__clkbuf_1
X_7314_ _3524_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__clkbuf_1
X_5575_ reg_data\[16\]\[18\] _1799_ _1800_ reg_data\[9\]\[18\] vssd1 vssd1 vccd1 vccd1
+ _2166_ sky130_fd_sc_hd__a22o_1
X_8294_ _4061_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__clkbuf_1
X_4526_ _1147_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__clkbuf_4
X_7245_ _3487_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__clkbuf_1
X_4457_ _1067_ _1079_ _1052_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__and3_2
X_7176_ reg_data\[7\]\[28\] _3187_ _3442_ vssd1 vssd1 vccd1 vccd1 _3451_ sky130_fd_sc_hd__mux2_1
X_6127_ reg_data\[16\]\[27\] _2405_ _2406_ reg_data\[9\]\[27\] vssd1 vssd1 vccd1 vccd1
+ _2700_ sky130_fd_sc_hd__a22o_1
X_4388_ _1015_ vssd1 vssd1 vccd1 vccd1 rs1_mux\[0\] sky130_fd_sc_hd__clkinv_2
X_6058_ reg_data\[30\]\[26\] _2204_ _1254_ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__and3_1
X_5009_ reg_data\[8\]\[9\] _1116_ _1119_ reg_data\[10\]\[9\] _1617_ vssd1 vssd1 vccd1
+ vccd1 _1618_ sky130_fd_sc_hd__a221o_1
X_9817_ clknet_leaf_51_i_clk rdata2\[1\] vssd1 vssd1 vccd1 vccd1 r_data2\[1\] sky130_fd_sc_hd__dfxtp_1
X_9748_ clknet_leaf_16_i_clk _0892_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_9679_ clknet_leaf_30_i_clk _0823_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_5360_ _1163_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__clkbuf_4
X_5291_ reg_data\[6\]\[13\] _1347_ _1632_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__and3_1
X_7030_ _3372_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__clkbuf_1
X_8981_ clknet_leaf_37_i_clk _0125_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_7932_ _3262_ reg_data\[28\]\[29\] _3844_ vssd1 vssd1 vccd1 vccd1 _3854_ sky130_fd_sc_hd__mux2_1
X_7863_ _3262_ reg_data\[27\]\[29\] _3807_ vssd1 vssd1 vccd1 vccd1 _3817_ sky130_fd_sc_hd__mux2_1
X_6814_ _3252_ reg_data\[22\]\[24\] _3244_ vssd1 vssd1 vccd1 vccd1 _3253_ sky130_fd_sc_hd__mux2_1
X_7794_ _3780_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__clkbuf_1
X_9602_ clknet_leaf_62_i_clk _0746_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6745_ i_data[2] vssd1 vssd1 vccd1 vccd1 _3206_ sky130_fd_sc_hd__clkbuf_4
X_9533_ clknet_leaf_4_i_clk _0677_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_9464_ clknet_leaf_10_i_clk _0608_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6676_ _3157_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__clkbuf_1
X_8415_ _3892_ reg_data\[17\]\[16\] _4119_ vssd1 vssd1 vccd1 vccd1 _4126_ sky130_fd_sc_hd__mux2_1
X_9395_ clknet_leaf_35_i_clk _0539_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5627_ reg_data\[7\]\[19\] _1780_ _2212_ _2213_ _2215_ vssd1 vssd1 vccd1 vccd1 _2216_
+ sky130_fd_sc_hd__a2111o_1
X_5558_ reg_data\[30\]\[18\] _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__and3_1
X_8346_ _4089_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__clkbuf_1
X_8277_ _4052_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__clkbuf_1
X_4509_ _1131_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__clkbuf_4
X_7228_ reg_data\[6\]\[20\] _3170_ _3478_ vssd1 vssd1 vccd1 vccd1 _3479_ sky130_fd_sc_hd__mux2_1
X_5489_ _2074_ _2078_ _2080_ _2082_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__or4_1
X_7159_ _3419_ vssd1 vssd1 vccd1 vccd1 _3442_ sky130_fd_sc_hd__buf_4
X_4860_ reg_data\[8\]\[6\] _1214_ _1217_ reg_data\[10\]\[6\] _1473_ vssd1 vssd1 vccd1
+ vccd1 _1474_ sky130_fd_sc_hd__a221o_1
X_6530_ r_data1\[20\] _3068_ vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__and2_1
X_4791_ _1160_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__clkbuf_4
X_6461_ reg_data\[25\]\[1\] _1140_ _3018_ _3019_ _3020_ vssd1 vssd1 vccd1 vccd1 _3021_
+ sky130_fd_sc_hd__a2111o_1
X_6392_ reg_data\[7\]\[0\] _1080_ _2952_ _2953_ _2954_ vssd1 vssd1 vccd1 vccd1 _2955_
+ sky130_fd_sc_hd__a2111o_1
X_5412_ reg_data\[20\]\[15\] _1629_ _1743_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__and3_1
X_8200_ _3882_ reg_data\[14\]\[11\] _4010_ vssd1 vssd1 vccd1 vccd1 _4012_ sky130_fd_sc_hd__mux2_1
X_9180_ clknet_leaf_5_i_clk _0324_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_5343_ _1941_ vssd1 vssd1 vccd1 vccd1 rdata1\[14\] sky130_fd_sc_hd__clkbuf_1
X_8131_ _3975_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__clkbuf_1
X_5274_ reg_data\[1\]\[13\] _1729_ _1793_ _1794_ reg_data\[15\]\[13\] vssd1 vssd1
+ vccd1 vccd1 _1875_ sky130_fd_sc_hd__a32o_1
X_8062_ _3938_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__clkbuf_1
X_7013_ _3363_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__clkbuf_1
X_8964_ clknet_leaf_62_i_clk _0108_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8895_ clknet_leaf_67_i_clk _0039_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_7915_ _3845_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__clkbuf_1
X_7846_ _3808_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__clkbuf_1
X_4989_ reg_data\[20\]\[9\] _1597_ _1315_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__and3_1
X_7777_ _3243_ reg_data\[26\]\[20\] _3771_ vssd1 vssd1 vccd1 vccd1 _3772_ sky130_fd_sc_hd__mux2_1
X_6728_ _3192_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__clkbuf_1
X_9516_ clknet_leaf_25_i_clk _0660_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_9447_ clknet_leaf_52_i_clk _0591_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6659_ reg_data\[4\]\[8\] _3145_ _3129_ vssd1 vssd1 vccd1 vccd1 _3146_ sky130_fd_sc_hd__mux2_1
X_9378_ clknet_leaf_60_i_clk _0522_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8329_ _4080_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__clkbuf_1
X_5961_ reg_data\[1\]\[24\] _2336_ _2399_ _2400_ reg_data\[15\]\[24\] vssd1 vssd1
+ vccd1 vccd1 _2540_ sky130_fd_sc_hd__a32o_1
X_8680_ _4266_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__clkbuf_1
X_7700_ _3235_ reg_data\[25\]\[16\] _3724_ vssd1 vssd1 vccd1 vccd1 _3731_ sky130_fd_sc_hd__mux2_1
X_4912_ reg_data\[12\]\[7\] _1354_ _1226_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__and3_1
X_5892_ _1071_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__buf_2
X_7631_ _3694_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__clkbuf_1
X_4843_ reg_data\[20\]\[6\] _1166_ _1180_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__and3_1
X_4774_ reg_data\[8\]\[5\] _1116_ _1119_ reg_data\[10\]\[5\] _1390_ vssd1 vssd1 vccd1
+ vccd1 _1391_ sky130_fd_sc_hd__a221o_1
X_7562_ _3657_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__clkbuf_1
X_9301_ clknet_leaf_35_i_clk _0445_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6513_ r_data1\[12\] _3057_ vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__and2_1
X_7493_ _3620_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__clkbuf_1
X_9232_ clknet_leaf_22_i_clk _0376_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6444_ reg_data\[12\]\[1\] _1082_ _1083_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__and3_1
X_6375_ _2930_ _2934_ _2936_ _2938_ vssd1 vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__or4_1
X_9163_ clknet_leaf_43_i_clk _0307_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5326_ _1043_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__buf_2
X_8114_ _3966_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__clkbuf_1
X_9094_ clknet_leaf_48_i_clk _0238_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8045_ _3929_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__clkbuf_1
X_5257_ reg_data\[18\]\[13\] _1656_ _1483_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__and3_1
X_5188_ _1105_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__clkbuf_4
X_8947_ clknet_leaf_36_i_clk _0091_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_8878_ clknet_leaf_29_i_clk _0022_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_7829_ _3799_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__clkbuf_1
X_4490_ reg_data\[27\]\[2\] _1096_ _1102_ _1107_ _1112_ vssd1 vssd1 vccd1 vccd1 _1113_
+ sky130_fd_sc_hd__a2111o_1
X_6160_ reg_data\[22\]\[28\] _1097_ _2256_ vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__and3_1
X_5111_ _1047_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__clkbuf_4
X_6091_ reg_data\[13\]\[26\] _2183_ _2299_ vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__and3_1
X_5042_ _1641_ _1645_ _1647_ _1649_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__or4_4
X_9850_ clknet_leaf_24_i_clk rs1_mux\[2\] vssd1 vssd1 vccd1 vccd1 rs1\[2\] sky130_fd_sc_hd__dfxtp_1
X_8801_ _4330_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__clkbuf_1
X_9781_ clknet_leaf_36_i_clk _0925_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6993_ reg_data\[0\]\[7\] _3143_ _3345_ vssd1 vssd1 vccd1 vccd1 _3353_ sky130_fd_sc_hd__mux2_1
X_5944_ reg_data\[18\]\[24\] _2261_ _2090_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__and3_1
X_8732_ _3869_ reg_data\[29\]\[5\] _4288_ vssd1 vssd1 vccd1 vccd1 _4294_ sky130_fd_sc_hd__mux2_1
X_5875_ reg_data\[26\]\[22\] _2455_ _2456_ reg_data\[29\]\[22\] vssd1 vssd1 vccd1
+ vccd1 _2457_ sky130_fd_sc_hd__a22o_1
X_8663_ _4257_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__clkbuf_1
X_7614_ _3685_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__clkbuf_1
X_4826_ _1428_ _1432_ _1436_ _1440_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__or4_1
X_8594_ _3867_ reg_data\[12\]\[4\] _4216_ vssd1 vssd1 vccd1 vccd1 _4221_ sky130_fd_sc_hd__mux2_1
X_7545_ _3648_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__clkbuf_1
X_4757_ reg_data\[3\]\[5\] _1054_ _1371_ _1372_ _1373_ vssd1 vssd1 vccd1 vccd1 _1374_
+ sky130_fd_sc_hd__a2111o_1
X_7476_ _3611_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__clkbuf_1
X_4688_ reg_data\[22\]\[4\] _1039_ _1236_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__and3_1
X_6427_ reg_data\[26\]\[0\] _1229_ _1231_ reg_data\[29\]\[0\] vssd1 vssd1 vccd1 vccd1
+ _2989_ sky130_fd_sc_hd__a22o_1
X_9215_ clknet_leaf_66_i_clk _0359_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6358_ reg_data\[6\]\[31\] _2555_ _1270_ vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__and3_1
X_9146_ clknet_leaf_10_i_clk _0290_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_5309_ reg_data\[8\]\[13\] _1841_ _1842_ reg_data\[10\]\[13\] _1908_ vssd1 vssd1
+ vccd1 vccd1 _1909_ sky130_fd_sc_hd__a221o_1
X_9077_ clknet_leaf_16_i_clk _0221_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6289_ reg_data\[16\]\[30\] _2405_ _2406_ reg_data\[9\]\[30\] vssd1 vssd1 vccd1 vccd1
+ _2856_ sky130_fd_sc_hd__a22o_1
X_8028_ _3918_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__clkbuf_1
X_5660_ reg_data\[2\]\[19\] _1837_ _1901_ _1902_ reg_data\[11\]\[19\] vssd1 vssd1
+ vccd1 vccd1 _2248_ sky130_fd_sc_hd__a32o_1
X_4611_ reg_data\[26\]\[2\] _1230_ _1232_ reg_data\[29\]\[2\] vssd1 vssd1 vccd1 vccd1
+ _1233_ sky130_fd_sc_hd__a22o_1
X_5591_ reg_data\[5\]\[18\] _1824_ _1954_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__and3_1
X_4542_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__buf_4
X_7330_ _3533_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__clkbuf_1
X_4473_ _1095_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__buf_4
X_7261_ reg_data\[5\]\[3\] _3135_ _3493_ vssd1 vssd1 vccd1 vccd1 _3497_ sky130_fd_sc_hd__mux2_1
X_6212_ _2773_ _2777_ _2779_ _2781_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__or4_1
X_9000_ clknet_leaf_49_i_clk _0144_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_7192_ reg_data\[6\]\[3\] _3135_ _3456_ vssd1 vssd1 vccd1 vccd1 _3460_ sky130_fd_sc_hd__mux2_1
X_6143_ reg_data\[5\]\[27\] _2430_ _1338_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__and3_1
X_6074_ reg_data\[8\]\[26\] _2403_ _2404_ reg_data\[10\]\[26\] _2648_ vssd1 vssd1
+ vccd1 vccd1 _2649_ sky130_fd_sc_hd__a221o_1
X_9902_ clknet_leaf_60_i_clk _0972_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_5025_ reg_data\[6\]\[9\] _1347_ _1632_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__and3_1
X_9833_ clknet_leaf_50_i_clk rdata2\[17\] vssd1 vssd1 vccd1 vccd1 r_data2\[17\] sky130_fd_sc_hd__dfxtp_1
X_6976_ _3343_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__clkbuf_1
X_9764_ clknet_leaf_60_i_clk _0908_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8715_ _4284_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__clkbuf_1
X_5927_ _1168_ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__buf_4
X_9695_ clknet_leaf_0_i_clk _0839_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8646_ _3919_ reg_data\[12\]\[29\] _4238_ vssd1 vssd1 vccd1 vccd1 _4248_ sky130_fd_sc_hd__mux2_1
X_5858_ _1205_ vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__buf_2
X_8577_ _4211_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__clkbuf_1
X_5789_ _1038_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__clkbuf_4
X_4809_ _1424_ vssd1 vssd1 vccd1 vccd1 rdata2\[5\] sky130_fd_sc_hd__clkbuf_1
X_7528_ _3198_ _3638_ vssd1 vssd1 vccd1 vccd1 _3639_ sky130_fd_sc_hd__and2_4
X_7459_ _3198_ _3601_ vssd1 vssd1 vccd1 vccd1 _3602_ sky130_fd_sc_hd__nand2_2
X_9129_ clknet_leaf_44_i_clk _0273_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_7__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_6830_ _3263_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__clkbuf_1
X_6761_ _3216_ reg_data\[22\]\[7\] _3202_ vssd1 vssd1 vccd1 vccd1 _3217_ sky130_fd_sc_hd__mux2_1
X_8500_ _3909_ reg_data\[18\]\[24\] _4166_ vssd1 vssd1 vccd1 vccd1 _4171_ sky130_fd_sc_hd__mux2_1
X_5712_ reg_data\[0\]\[20\] _1821_ _2295_ _2296_ _2297_ vssd1 vssd1 vccd1 vccd1 _2298_
+ sky130_fd_sc_hd__a2111o_1
X_6692_ i_data[19] vssd1 vssd1 vccd1 vccd1 _3168_ sky130_fd_sc_hd__clkbuf_4
X_9480_ clknet_leaf_46_i_clk _0624_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_8431_ _4134_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__clkbuf_1
X_5643_ reg_data\[25\]\[19\] _1810_ _2228_ _2229_ _2230_ vssd1 vssd1 vccd1 vccd1 _2231_
+ sky130_fd_sc_hd__a2111o_1
X_8362_ _3907_ reg_data\[16\]\[23\] _4094_ vssd1 vssd1 vccd1 vccd1 _4098_ sky130_fd_sc_hd__mux2_1
X_5574_ reg_data\[27\]\[18\] _1786_ _2162_ _2163_ _2164_ vssd1 vssd1 vccd1 vccd1 _2165_
+ sky130_fd_sc_hd__a2111o_1
X_7313_ reg_data\[5\]\[28\] _3187_ _3515_ vssd1 vssd1 vccd1 vccd1 _3524_ sky130_fd_sc_hd__mux2_1
X_4525_ rs2_mux\[0\] _1005_ _1010_ _1013_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__and4_2
X_8293_ _3907_ reg_data\[15\]\[23\] _4057_ vssd1 vssd1 vccd1 vccd1 _4061_ sky130_fd_sc_hd__mux2_1
X_7244_ reg_data\[6\]\[28\] _3187_ _3478_ vssd1 vssd1 vccd1 vccd1 _3487_ sky130_fd_sc_hd__mux2_1
X_4456_ _1030_ rs1_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__nor2_1
X_7175_ _3450_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__clkbuf_1
X_4387_ _1014_ i_rs1[0] i_rs_valid vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__mux2_2
X_6126_ reg_data\[27\]\[27\] _2392_ _2696_ _2697_ _2698_ vssd1 vssd1 vccd1 vccd1 _2699_
+ sky130_fd_sc_hd__a2111o_1
X_6057_ reg_data\[20\]\[26\] _2524_ _1059_ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__and3_1
X_5008_ reg_data\[16\]\[9\] _1121_ _1123_ reg_data\[9\]\[9\] vssd1 vssd1 vccd1 vccd1
+ _1617_ sky130_fd_sc_hd__a22o_1
X_9816_ clknet_leaf_50_i_clk rdata2\[0\] vssd1 vssd1 vccd1 vccd1 r_data2\[0\] sky130_fd_sc_hd__dfxtp_1
X_9747_ clknet_leaf_17_i_clk _0891_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6959_ _3250_ reg_data\[10\]\[23\] _3331_ vssd1 vssd1 vccd1 vccd1 _3335_ sky130_fd_sc_hd__mux2_1
X_9678_ clknet_leaf_30_i_clk _0822_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_8629_ _4239_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_31_i_clk clknet_3_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_46_i_clk clknet_3_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5290_ reg_data\[3\]\[13\] _1815_ _1887_ _1888_ _1889_ vssd1 vssd1 vccd1 vccd1 _1890_
+ sky130_fd_sc_hd__a2111o_1
X_8980_ clknet_leaf_32_i_clk _0124_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_7931_ _3853_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__clkbuf_1
X_7862_ _3816_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__clkbuf_1
X_9601_ clknet_leaf_73_i_clk _0745_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_7793_ _3260_ reg_data\[26\]\[28\] _3771_ vssd1 vssd1 vccd1 vccd1 _3780_ sky130_fd_sc_hd__mux2_1
X_6813_ i_data[24] vssd1 vssd1 vccd1 vccd1 _3252_ sky130_fd_sc_hd__buf_2
X_6744_ _3205_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__clkbuf_1
X_9532_ clknet_leaf_11_i_clk _0676_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_9463_ clknet_leaf_43_i_clk _0607_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6675_ reg_data\[4\]\[13\] _3156_ _3150_ vssd1 vssd1 vccd1 vccd1 _3157_ sky130_fd_sc_hd__mux2_1
X_5626_ reg_data\[13\]\[19\] _2214_ _2102_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__and3_1
X_8414_ _4125_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__clkbuf_1
X_9394_ clknet_leaf_33_i_clk _0538_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_5557_ reg_data\[18\]\[18\] _1656_ _2090_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__and3_1
X_8345_ _3890_ reg_data\[16\]\[15\] _4083_ vssd1 vssd1 vccd1 vccd1 _4089_ sky130_fd_sc_hd__mux2_1
X_4508_ _1097_ _1117_ _1094_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__and3_4
X_8276_ _3890_ reg_data\[15\]\[15\] _4046_ vssd1 vssd1 vccd1 vccd1 _4052_ sky130_fd_sc_hd__mux2_1
X_5488_ reg_data\[24\]\[16\] _1847_ _1848_ reg_data\[28\]\[16\] _2081_ vssd1 vssd1
+ vccd1 vccd1 _2082_ sky130_fd_sc_hd__a221o_1
X_7227_ _3455_ vssd1 vssd1 vccd1 vccd1 _3478_ sky130_fd_sc_hd__buf_4
X_4439_ _1034_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__clkbuf_4
X_7158_ _3441_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__clkbuf_1
X_6109_ reg_data\[25\]\[27\] _2370_ _2679_ _2680_ _2681_ vssd1 vssd1 vccd1 vccd1 _2682_
+ sky130_fd_sc_hd__a2111o_1
X_7089_ _3404_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__clkbuf_1
X_4790_ reg_data\[6\]\[5\] _1347_ _1152_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__and3_1
X_6460_ reg_data\[17\]\[1\] _1162_ _1148_ vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__and3_1
X_6391_ reg_data\[13\]\[0\] _1076_ _1087_ vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__and3_1
X_5411_ reg_data\[30\]\[15\] _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__and3_1
X_5342_ _1932_ _1936_ _1938_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__or4_1
X_8130_ _3879_ reg_data\[13\]\[10\] _3974_ vssd1 vssd1 vccd1 vccd1 _3975_ sky130_fd_sc_hd__mux2_1
X_8061_ _3879_ reg_data\[30\]\[10\] _3937_ vssd1 vssd1 vccd1 vccd1 _3938_ sky130_fd_sc_hd__mux2_1
X_5273_ reg_data\[2\]\[13\] _1613_ _1790_ _1791_ reg_data\[11\]\[13\] vssd1 vssd1
+ vccd1 vccd1 _1874_ sky130_fd_sc_hd__a32o_1
X_7012_ reg_data\[0\]\[16\] _3162_ _3356_ vssd1 vssd1 vccd1 vccd1 _3363_ sky130_fd_sc_hd__mux2_1
X_8963_ clknet_leaf_59_i_clk _0107_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8894_ clknet_leaf_6_i_clk _0038_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_7914_ _3243_ reg_data\[28\]\[20\] _3844_ vssd1 vssd1 vccd1 vccd1 _3845_ sky130_fd_sc_hd__mux2_1
X_7845_ _3243_ reg_data\[27\]\[20\] _3807_ vssd1 vssd1 vccd1 vccd1 _3808_ sky130_fd_sc_hd__mux2_1
X_9515_ clknet_leaf_25_i_clk _0659_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_7776_ _3748_ vssd1 vssd1 vccd1 vccd1 _3771_ sky130_fd_sc_hd__buf_4
X_4988_ _1034_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__buf_2
X_6727_ reg_data\[4\]\[30\] _3191_ _3128_ vssd1 vssd1 vccd1 vccd1 _3192_ sky130_fd_sc_hd__mux2_1
X_6658_ i_data[8] vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__clkbuf_4
X_9446_ clknet_leaf_51_i_clk _0590_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_5609_ reg_data\[22\]\[19\] _2143_ _1651_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__and3_1
X_9377_ clknet_leaf_1_i_clk _0521_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6589_ _3100_ vssd1 vssd1 vccd1 vccd1 o_data2[15] sky130_fd_sc_hd__buf_2
X_8328_ _3873_ reg_data\[16\]\[7\] _4072_ vssd1 vssd1 vccd1 vccd1 _4080_ sky130_fd_sc_hd__mux2_1
X_8259_ _3873_ reg_data\[15\]\[7\] _4035_ vssd1 vssd1 vccd1 vccd1 _4043_ sky130_fd_sc_hd__mux2_1
X_5960_ reg_data\[2\]\[24\] _2219_ _2396_ _2397_ reg_data\[11\]\[24\] vssd1 vssd1
+ vccd1 vccd1 _2539_ sky130_fd_sc_hd__a32o_1
X_5891_ reg_data\[0\]\[23\] _2381_ _2468_ _2470_ _2471_ vssd1 vssd1 vccd1 vccd1 _2472_
+ sky130_fd_sc_hd__a2111o_1
X_4911_ reg_data\[14\]\[7\] _1189_ _1193_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__and3_1
X_7630_ _3233_ reg_data\[24\]\[15\] _3688_ vssd1 vssd1 vccd1 vccd1 _3694_ sky130_fd_sc_hd__mux2_1
X_4842_ reg_data\[30\]\[6\] _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__and3_1
X_4773_ reg_data\[16\]\[5\] _1121_ _1123_ reg_data\[9\]\[5\] vssd1 vssd1 vccd1 vccd1
+ _1390_ sky130_fd_sc_hd__a22o_1
X_7561_ reg_data\[23\]\[15\] _3160_ _3651_ vssd1 vssd1 vccd1 vccd1 _3657_ sky130_fd_sc_hd__mux2_1
X_9300_ clknet_leaf_33_i_clk _0444_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6512_ _3059_ vssd1 vssd1 vccd1 vccd1 o_data1[11] sky130_fd_sc_hd__buf_2
X_7492_ _3233_ reg_data\[21\]\[15\] _3614_ vssd1 vssd1 vccd1 vccd1 _3620_ sky130_fd_sc_hd__mux2_1
X_9231_ clknet_leaf_30_i_clk _0375_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6443_ reg_data\[14\]\[1\] _1074_ _1313_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__and3_1
X_6374_ reg_data\[24\]\[31\] _2453_ _2454_ reg_data\[28\]\[31\] _2937_ vssd1 vssd1
+ vccd1 vccd1 _2938_ sky130_fd_sc_hd__a221o_1
X_9162_ clknet_leaf_43_i_clk _0306_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8113_ _3863_ reg_data\[13\]\[2\] _3963_ vssd1 vssd1 vccd1 vccd1 _3966_ sky130_fd_sc_hd__mux2_1
X_9093_ clknet_leaf_62_i_clk _0237_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5325_ reg_data\[4\]\[14\] _1718_ _1863_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__and3_1
X_5256_ reg_data\[25\]\[13\] _1764_ _1854_ _1855_ _1856_ vssd1 vssd1 vccd1 vccd1 _1857_
+ sky130_fd_sc_hd__a2111o_1
X_8044_ _3863_ reg_data\[30\]\[2\] _3926_ vssd1 vssd1 vccd1 vccd1 _3929_ sky130_fd_sc_hd__mux2_1
X_5187_ _1064_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__clkbuf_4
X_8946_ clknet_leaf_36_i_clk _0090_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_8877_ clknet_leaf_25_i_clk _0021_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_7828_ _3227_ reg_data\[27\]\[12\] _3796_ vssd1 vssd1 vccd1 vccd1 _3799_ sky130_fd_sc_hd__mux2_1
X_7759_ _3762_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__clkbuf_1
X_9429_ clknet_leaf_34_i_clk _0573_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6090_ reg_data\[0\]\[26\] _2427_ _2661_ _2662_ _2663_ vssd1 vssd1 vccd1 vccd1 _2664_
+ sky130_fd_sc_hd__a2111o_1
X_5110_ reg_data\[3\]\[11\] _1054_ _1712_ _1713_ _1714_ vssd1 vssd1 vccd1 vccd1 _1715_
+ sky130_fd_sc_hd__a2111o_1
X_5041_ reg_data\[24\]\[9\] _1225_ _1228_ reg_data\[28\]\[9\] _1648_ vssd1 vssd1 vccd1
+ vccd1 _1649_ sky130_fd_sc_hd__a221o_1
X_9780_ clknet_leaf_37_i_clk _0924_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_8800_ reg_data\[11\]\[5\] i_data[5] _4324_ vssd1 vssd1 vccd1 vccd1 _4330_ sky130_fd_sc_hd__mux2_1
X_8731_ _4293_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__clkbuf_1
X_6992_ _3352_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__clkbuf_1
X_5943_ reg_data\[25\]\[24\] _2370_ _2519_ _2520_ _2521_ vssd1 vssd1 vccd1 vccd1 _2522_
+ sky130_fd_sc_hd__a2111o_1
X_5874_ _1231_ vssd1 vssd1 vccd1 vccd1 _2456_ sky130_fd_sc_hd__clkbuf_4
X_8662_ reg_data\[19\]\[4\] _3137_ _4252_ vssd1 vssd1 vccd1 vccd1 _4257_ sky130_fd_sc_hd__mux2_1
X_7613_ _3216_ reg_data\[24\]\[7\] _3677_ vssd1 vssd1 vccd1 vccd1 _3685_ sky130_fd_sc_hd__mux2_1
X_4825_ reg_data\[7\]\[6\] _1081_ _1437_ _1438_ _1439_ vssd1 vssd1 vccd1 vccd1 _1440_
+ sky130_fd_sc_hd__a2111o_1
X_8593_ _4220_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__clkbuf_1
X_7544_ reg_data\[23\]\[7\] _3143_ _3640_ vssd1 vssd1 vccd1 vccd1 _3648_ sky130_fd_sc_hd__mux2_1
X_4756_ reg_data\[30\]\[5\] _1062_ _1090_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__and3_1
X_4687_ _1306_ vssd1 vssd1 vccd1 vccd1 rdata2\[3\] sky130_fd_sc_hd__clkbuf_1
X_7475_ _3216_ reg_data\[21\]\[7\] _3603_ vssd1 vssd1 vccd1 vccd1 _3611_ sky130_fd_sc_hd__mux2_1
X_6426_ reg_data\[8\]\[0\] _1213_ _1216_ reg_data\[10\]\[0\] _2987_ vssd1 vssd1 vccd1
+ vccd1 _2988_ sky130_fd_sc_hd__a221o_1
X_9214_ clknet_leaf_6_i_clk _0358_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6357_ reg_data\[3\]\[31\] _2421_ _2918_ _2919_ _2920_ vssd1 vssd1 vccd1 vccd1 _2921_
+ sky130_fd_sc_hd__a2111o_1
X_9145_ clknet_leaf_11_i_clk _0289_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_5308_ reg_data\[16\]\[13\] _1843_ _1844_ reg_data\[9\]\[13\] vssd1 vssd1 vccd1 vccd1
+ _1908_ sky130_fd_sc_hd__a22o_1
X_9076_ clknet_leaf_16_i_clk _0220_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6288_ reg_data\[27\]\[30\] _2392_ _2852_ _2853_ _2854_ vssd1 vssd1 vccd1 vccd1 _2855_
+ sky130_fd_sc_hd__a2111o_1
X_8027_ _3917_ reg_data\[9\]\[28\] _3901_ vssd1 vssd1 vccd1 vccd1 _3918_ sky130_fd_sc_hd__mux2_1
X_5239_ _1213_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__clkbuf_4
X_8929_ clknet_leaf_1_i_clk _0073_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_4610_ _1231_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__clkbuf_4
X_5590_ reg_data\[4\]\[18\] _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__and3_1
X_4541_ rs2_mux\[0\] _1005_ rs2_mux\[2\] rs2_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1163_
+ sky130_fd_sc_hd__and4bb_4
X_4472_ _1062_ _1094_ _1052_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__and3_4
X_7260_ _3496_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__clkbuf_1
X_6211_ reg_data\[24\]\[28\] _2453_ _2454_ reg_data\[28\]\[28\] _2780_ vssd1 vssd1
+ vccd1 vccd1 _2781_ sky130_fd_sc_hd__a221o_1
X_7191_ _3459_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__clkbuf_1
X_6142_ reg_data\[4\]\[27\] _1175_ _1342_ vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__and3_1
X_6073_ reg_data\[16\]\[26\] _2405_ _2406_ reg_data\[9\]\[26\] vssd1 vssd1 vccd1 vccd1
+ _2648_ sky130_fd_sc_hd__a22o_1
X_5024_ _1151_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__clkbuf_4
X_9901_ clknet_leaf_61_i_clk _0971_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_9832_ clknet_leaf_50_i_clk rdata2\[16\] vssd1 vssd1 vccd1 vccd1 r_data2\[16\] sky130_fd_sc_hd__dfxtp_1
X_6975_ _3266_ reg_data\[10\]\[31\] _3308_ vssd1 vssd1 vccd1 vccd1 _3343_ sky130_fd_sc_hd__mux2_1
X_9763_ clknet_leaf_60_i_clk _0907_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_5926_ reg_data\[23\]\[23\] _2440_ _2441_ reg_data\[19\]\[23\] vssd1 vssd1 vccd1
+ vccd1 _2506_ sky130_fd_sc_hd__a22o_1
X_8714_ reg_data\[19\]\[29\] _3189_ _4274_ vssd1 vssd1 vccd1 vccd1 _4284_ sky130_fd_sc_hd__mux2_1
X_9694_ clknet_leaf_76_i_clk _0838_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8645_ _4247_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__clkbuf_1
X_5857_ _1198_ vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__clkbuf_4
X_8576_ reg_data\[1\]\[28\] _3187_ _4202_ vssd1 vssd1 vccd1 vccd1 _4211_ sky130_fd_sc_hd__mux2_1
X_5788_ reg_data\[22\]\[22\] _2143_ _2256_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__and3_1
X_4808_ _1415_ _1419_ _1421_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__or4_1
X_7527_ i_rd[0] i_rd[1] _3126_ vssd1 vssd1 vccd1 vccd1 _3638_ sky130_fd_sc_hd__nor3_4
X_4739_ _1340_ _1346_ _1351_ _1356_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__or4_1
X_7458_ _3600_ vssd1 vssd1 vccd1 vccd1 _3601_ sky130_fd_sc_hd__buf_2
X_6409_ reg_data\[30\]\[0\] _1146_ _1163_ vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__and3_1
X_7389_ _3381_ _3198_ vssd1 vssd1 vccd1 vccd1 _3564_ sky130_fd_sc_hd__nand2_4
X_9128_ clknet_leaf_46_i_clk _0272_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_9059_ clknet_leaf_66_i_clk _0203_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6760_ i_data[7] vssd1 vssd1 vccd1 vccd1 _3216_ sky130_fd_sc_hd__buf_2
X_5711_ reg_data\[5\]\[20\] _1824_ _1954_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__and3_1
X_6691_ _3167_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__clkbuf_1
X_8430_ _3907_ reg_data\[17\]\[23\] _4130_ vssd1 vssd1 vccd1 vccd1 _4134_ sky130_fd_sc_hd__mux2_1
X_5642_ reg_data\[17\]\[19\] _2117_ _1275_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__and3_1
X_8361_ _4097_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__clkbuf_1
X_5573_ reg_data\[1\]\[18\] _1729_ _1793_ _1794_ reg_data\[15\]\[18\] vssd1 vssd1
+ vccd1 vccd1 _2164_ sky130_fd_sc_hd__a32o_1
X_7312_ _3523_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__clkbuf_1
X_4524_ _1142_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__buf_2
X_8292_ _4060_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__clkbuf_1
X_7243_ _3486_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__clkbuf_1
X_4455_ reg_data\[0\]\[2\] _1070_ _1073_ _1075_ _1077_ vssd1 vssd1 vccd1 vccd1 _1078_
+ sky130_fd_sc_hd__a2111o_1
X_7174_ reg_data\[7\]\[27\] _3185_ _3442_ vssd1 vssd1 vccd1 vccd1 _3450_ sky130_fd_sc_hd__mux2_1
X_4386_ rs1\[0\] vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__clkinv_2
X_6125_ reg_data\[1\]\[27\] _2336_ _2399_ _2400_ reg_data\[15\]\[27\] vssd1 vssd1
+ vccd1 vccd1 _2698_ sky130_fd_sc_hd__a32o_1
X_6056_ reg_data\[18\]\[26\] _2261_ _2090_ vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__and3_1
X_5007_ reg_data\[27\]\[9\] _1096_ _1612_ _1614_ _1615_ vssd1 vssd1 vccd1 vccd1 _1616_
+ sky130_fd_sc_hd__a2111o_1
X_9815_ clknet_leaf_39_i_clk rdata1\[31\] vssd1 vssd1 vccd1 vccd1 r_data1\[31\] sky130_fd_sc_hd__dfxtp_1
X_9746_ clknet_leaf_17_i_clk _0890_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6958_ _3334_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__clkbuf_1
X_9677_ clknet_leaf_29_i_clk _0821_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6889_ reg_data\[2\]\[23\] _3177_ _3293_ vssd1 vssd1 vccd1 vccd1 _3297_ sky130_fd_sc_hd__mux2_1
X_5909_ _1142_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__clkbuf_4
X_8628_ _3900_ reg_data\[12\]\[20\] _4238_ vssd1 vssd1 vccd1 vccd1 _4239_ sky130_fd_sc_hd__mux2_1
X_8559_ _4179_ vssd1 vssd1 vccd1 vccd1 _4202_ sky130_fd_sc_hd__clkbuf_4
X_7930_ _3260_ reg_data\[28\]\[28\] _3844_ vssd1 vssd1 vccd1 vccd1 _3853_ sky130_fd_sc_hd__mux2_1
X_7861_ _3260_ reg_data\[27\]\[28\] _3807_ vssd1 vssd1 vccd1 vccd1 _3816_ sky130_fd_sc_hd__mux2_1
X_6812_ _3251_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__clkbuf_1
X_9600_ clknet_leaf_74_i_clk _0744_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7792_ _3779_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__clkbuf_1
X_9531_ clknet_leaf_4_i_clk _0675_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6743_ _3204_ reg_data\[22\]\[1\] _3202_ vssd1 vssd1 vccd1 vccd1 _3205_ sky130_fd_sc_hd__mux2_1
X_9462_ clknet_leaf_43_i_clk _0606_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6674_ i_data[13] vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__buf_2
X_5625_ _1067_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__clkbuf_4
X_8413_ _3890_ reg_data\[17\]\[15\] _4119_ vssd1 vssd1 vccd1 vccd1 _4125_ sky130_fd_sc_hd__mux2_1
X_9393_ clknet_leaf_35_i_clk _0537_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_5556_ reg_data\[25\]\[18\] _1764_ _2144_ _2145_ _2146_ vssd1 vssd1 vccd1 vccd1 _2147_
+ sky130_fd_sc_hd__a2111o_1
X_8344_ _4088_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__clkbuf_1
X_8275_ _4051_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__clkbuf_1
X_4507_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__clkbuf_4
X_5487_ reg_data\[26\]\[16\] _1849_ _1850_ reg_data\[29\]\[16\] vssd1 vssd1 vccd1
+ vccd1 _2081_ sky130_fd_sc_hd__a22o_1
X_7226_ _3477_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
X_4438_ reg_data\[20\]\[2\] _1058_ _1060_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__and3_1
X_4369_ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__buf_6
X_7157_ reg_data\[7\]\[19\] _3168_ _3431_ vssd1 vssd1 vccd1 vccd1 _3441_ sky130_fd_sc_hd__mux2_1
X_6108_ reg_data\[21\]\[27\] _1058_ _2087_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__and3_1
X_7088_ _3241_ reg_data\[8\]\[19\] _3394_ vssd1 vssd1 vccd1 vccd1 _3404_ sky130_fd_sc_hd__mux2_1
X_6039_ reg_data\[12\]\[25\] _2562_ _2016_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__and3_1
X_9729_ clknet_leaf_5_i_clk _0873_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6390_ reg_data\[12\]\[0\] _1082_ _1083_ vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__and3_1
X_5410_ _1163_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__buf_4
X_5341_ reg_data\[24\]\[14\] _1803_ _1804_ reg_data\[28\]\[14\] _1939_ vssd1 vssd1
+ vccd1 vccd1 _1940_ sky130_fd_sc_hd__a221o_1
X_8060_ _3925_ vssd1 vssd1 vccd1 vccd1 _3937_ sky130_fd_sc_hd__buf_4
X_5272_ reg_data\[23\]\[13\] _1787_ _1788_ reg_data\[19\]\[13\] vssd1 vssd1 vccd1
+ vccd1 _1873_ sky130_fd_sc_hd__a22o_1
X_7011_ _3362_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__clkbuf_1
X_8962_ clknet_leaf_62_i_clk _0106_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_7913_ _3821_ vssd1 vssd1 vccd1 vccd1 _3844_ sky130_fd_sc_hd__buf_4
X_8893_ clknet_leaf_67_i_clk _0037_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_30_i_clk clknet_3_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_7844_ _3784_ vssd1 vssd1 vccd1 vccd1 _3807_ sky130_fd_sc_hd__buf_4
X_7775_ _3770_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__clkbuf_1
X_6726_ i_data[30] vssd1 vssd1 vccd1 vccd1 _3191_ sky130_fd_sc_hd__buf_4
X_9514_ clknet_leaf_26_i_clk _0658_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_4987_ reg_data\[30\]\[9\] _1312_ _1313_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__and3_1
X_6657_ _3144_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__clkbuf_1
X_9445_ clknet_leaf_51_i_clk _0589_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_45_i_clk clknet_3_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_9376_ clknet_leaf_74_i_clk _0520_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_5608_ _2197_ vssd1 vssd1 vccd1 vccd1 rdata2\[18\] sky130_fd_sc_hd__clkbuf_1
X_6588_ r_data2\[15\] _3094_ vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__and2_1
X_8327_ _4079_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__clkbuf_1
X_5539_ reg_data\[12\]\[17\] _1960_ _2016_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__and3_1
X_8258_ _4042_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__clkbuf_1
X_7209_ reg_data\[6\]\[11\] _3152_ _3467_ vssd1 vssd1 vccd1 vccd1 _3469_ sky130_fd_sc_hd__mux2_1
X_8189_ _3871_ reg_data\[14\]\[6\] _3999_ vssd1 vssd1 vccd1 vccd1 _4006_ sky130_fd_sc_hd__mux2_1
X_5890_ reg_data\[5\]\[23\] _2097_ _1925_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__and3_1
X_4910_ reg_data\[13\]\[7\] _1186_ _1191_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__and3_1
X_4841_ reg_data\[18\]\[6\] _1159_ _1168_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__and3_1
X_7560_ _3656_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__clkbuf_1
X_4772_ reg_data\[27\]\[5\] _1096_ _1386_ _1387_ _1388_ vssd1 vssd1 vccd1 vccd1 _1389_
+ sky130_fd_sc_hd__a2111o_1
X_6511_ r_data1\[11\] _3057_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__and2_1
X_7491_ _3619_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__clkbuf_1
X_9230_ clknet_leaf_32_i_clk _0374_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6442_ reg_data\[0\]\[1\] _1069_ _3000_ _3001_ _3002_ vssd1 vssd1 vccd1 vccd1 _3003_
+ sky130_fd_sc_hd__a2111o_1
X_9161_ clknet_leaf_44_i_clk _0305_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6373_ reg_data\[26\]\[31\] _2455_ _2456_ reg_data\[29\]\[31\] vssd1 vssd1 vccd1
+ vccd1 _2937_ sky130_fd_sc_hd__a22o_1
X_8112_ _3965_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__clkbuf_1
X_9092_ clknet_leaf_62_i_clk _0236_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_5324_ reg_data\[6\]\[14\] _1600_ _1716_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__and3_1
X_8043_ _3928_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__clkbuf_1
X_5255_ reg_data\[17\]\[13\] _1480_ _1108_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__and3_1
X_5186_ reg_data\[23\]\[12\] _1787_ _1788_ reg_data\[19\]\[12\] vssd1 vssd1 vccd1
+ vccd1 _1789_ sky130_fd_sc_hd__a22o_1
X_8945_ clknet_leaf_36_i_clk _0089_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_8876_ clknet_leaf_27_i_clk _0020_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_7827_ _3798_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__clkbuf_1
X_7758_ _3225_ reg_data\[26\]\[11\] _3760_ vssd1 vssd1 vccd1 vccd1 _3762_ sky130_fd_sc_hd__mux2_1
X_6709_ reg_data\[4\]\[24\] _3179_ _3171_ vssd1 vssd1 vccd1 vccd1 _3180_ sky130_fd_sc_hd__mux2_1
X_7689_ _3725_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__clkbuf_1
X_9428_ clknet_leaf_31_i_clk _0572_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_9359_ clknet_leaf_31_i_clk _0503_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_5040_ reg_data\[26\]\[9\] _1230_ _1232_ reg_data\[29\]\[9\] vssd1 vssd1 vccd1 vccd1
+ _1648_ sky130_fd_sc_hd__a22o_1
X_6991_ reg_data\[0\]\[6\] _3141_ _3345_ vssd1 vssd1 vccd1 vccd1 _3352_ sky130_fd_sc_hd__mux2_1
X_5942_ reg_data\[21\]\[24\] _2086_ _2087_ vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__and3_1
X_8730_ _3867_ reg_data\[29\]\[4\] _4288_ vssd1 vssd1 vccd1 vccd1 _4293_ sky130_fd_sc_hd__mux2_1
X_5873_ _1229_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__clkbuf_4
X_8661_ _4256_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__clkbuf_1
X_7612_ _3684_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__clkbuf_1
X_4824_ reg_data\[13\]\[6\] _1089_ _1257_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__and3_1
X_8592_ _3865_ reg_data\[12\]\[3\] _4216_ vssd1 vssd1 vccd1 vccd1 _4220_ sky130_fd_sc_hd__mux2_1
X_7543_ _3647_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__clkbuf_1
X_4755_ reg_data\[20\]\[5\] _1312_ _1060_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__and3_1
X_4686_ _1293_ _1301_ _1303_ _1305_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__or4_2
X_7474_ _3610_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__clkbuf_1
X_9213_ clknet_leaf_67_i_clk _0357_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6425_ reg_data\[16\]\[0\] _1218_ _1220_ reg_data\[9\]\[0\] vssd1 vssd1 vccd1 vccd1
+ _2987_ sky130_fd_sc_hd__a22o_1
X_6356_ reg_data\[20\]\[31\] _1150_ _1283_ vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__and3_1
X_9144_ clknet_leaf_12_i_clk _0288_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_9075_ clknet_leaf_18_i_clk _0219_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5307_ reg_data\[27\]\[13\] _1833_ _1900_ _1903_ _1906_ vssd1 vssd1 vccd1 vccd1 _1907_
+ sky130_fd_sc_hd__a2111o_1
X_8026_ i_data[28] vssd1 vssd1 vccd1 vccd1 _3917_ sky130_fd_sc_hd__clkbuf_4
X_6287_ reg_data\[1\]\[30\] _2336_ _2399_ _2400_ reg_data\[15\]\[30\] vssd1 vssd1
+ vccd1 vccd1 _2854_ sky130_fd_sc_hd__a32o_1
X_5238_ reg_data\[27\]\[12\] _1833_ _1836_ _1838_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_
+ sky130_fd_sc_hd__a2111o_1
X_5169_ reg_data\[20\]\[12\] _1312_ _1060_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__and3_1
X_8928_ clknet_leaf_75_i_clk _0072_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8859_ clknet_leaf_0_i_clk _0003_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_4540_ _1138_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__buf_2
X_4471_ rs1_mux\[2\] _1033_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__nor2_2
X_6210_ reg_data\[26\]\[28\] _2455_ _2456_ reg_data\[29\]\[28\] vssd1 vssd1 vccd1
+ vccd1 _2780_ sky130_fd_sc_hd__a22o_1
X_7190_ reg_data\[6\]\[2\] _3133_ _3456_ vssd1 vssd1 vccd1 vccd1 _3459_ sky130_fd_sc_hd__mux2_1
X_6141_ reg_data\[6\]\[27\] _2555_ _2237_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__and3_1
X_6072_ reg_data\[27\]\[26\] _2392_ _2644_ _2645_ _2646_ vssd1 vssd1 vccd1 vccd1 _2647_
+ sky130_fd_sc_hd__a2111o_1
X_9900_ clknet_leaf_61_i_clk _0970_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_5023_ reg_data\[3\]\[9\] _1158_ _1627_ _1628_ _1630_ vssd1 vssd1 vccd1 vccd1 _1631_
+ sky130_fd_sc_hd__a2111o_1
X_9831_ clknet_leaf_50_i_clk rdata2\[15\] vssd1 vssd1 vccd1 vccd1 r_data2\[15\] sky130_fd_sc_hd__dfxtp_1
X_6974_ _3342_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__clkbuf_1
X_9762_ clknet_leaf_60_i_clk _0906_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_5925_ _2492_ _2496_ _2500_ _2504_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__or4_1
X_8713_ _4283_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__clkbuf_1
X_9693_ clknet_leaf_0_i_clk _0837_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_8644_ _3917_ reg_data\[12\]\[28\] _4238_ vssd1 vssd1 vccd1 vccd1 _4247_ sky130_fd_sc_hd__mux2_1
X_5856_ _2420_ _2426_ _2432_ _2437_ vssd1 vssd1 vccd1 vccd1 _2438_ sky130_fd_sc_hd__or4_2
X_4807_ reg_data\[24\]\[5\] _1225_ _1228_ reg_data\[28\]\[5\] _1422_ vssd1 vssd1 vccd1
+ vccd1 _1423_ sky130_fd_sc_hd__a221o_1
X_8575_ _4210_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__clkbuf_1
X_5787_ _1036_ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__clkbuf_4
X_7526_ _3637_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__clkbuf_1
X_4738_ reg_data\[7\]\[4\] _1185_ _1352_ _1353_ _1355_ vssd1 vssd1 vccd1 vccd1 _1356_
+ sky130_fd_sc_hd__a2111o_1
X_4669_ _1187_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__clkbuf_4
X_7457_ i_rd[0] i_rd[1] i_write i_reset_n vssd1 vssd1 vccd1 vccd1 _3600_ sky130_fd_sc_hd__and4b_1
X_6408_ reg_data\[18\]\[0\] _1143_ _1167_ vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__and3_1
X_7388_ _3563_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__clkbuf_1
X_9127_ clknet_leaf_46_i_clk _0271_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6339_ reg_data\[23\]\[31\] _2393_ _2394_ reg_data\[19\]\[31\] vssd1 vssd1 vccd1
+ vccd1 _2904_ sky130_fd_sc_hd__a22o_1
X_9058_ clknet_leaf_66_i_clk _0202_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8009_ _3905_ reg_data\[9\]\[22\] _3901_ vssd1 vssd1 vccd1 vccd1 _3906_ sky130_fd_sc_hd__mux2_1
X_5710_ reg_data\[4\]\[20\] _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__and3_1
X_6690_ reg_data\[4\]\[18\] _3166_ _3150_ vssd1 vssd1 vccd1 vccd1 _3167_ sky130_fd_sc_hd__mux2_1
X_5641_ reg_data\[21\]\[19\] _1883_ _1943_ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__and3_1
X_8360_ _3905_ reg_data\[16\]\[22\] _4094_ vssd1 vssd1 vccd1 vccd1 _4097_ sky130_fd_sc_hd__mux2_1
X_5572_ reg_data\[2\]\[18\] _1613_ _1790_ _1791_ reg_data\[11\]\[18\] vssd1 vssd1
+ vccd1 vccd1 _2163_ sky130_fd_sc_hd__a32o_1
X_7311_ reg_data\[5\]\[27\] _3185_ _3515_ vssd1 vssd1 vccd1 vccd1 _3523_ sky130_fd_sc_hd__mux2_1
X_8291_ _3905_ reg_data\[15\]\[22\] _4057_ vssd1 vssd1 vccd1 vccd1 _4060_ sky130_fd_sc_hd__mux2_1
X_4523_ reg_data\[21\]\[2\] _1143_ _1144_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__and3_1
X_7242_ reg_data\[6\]\[27\] _3185_ _3478_ vssd1 vssd1 vccd1 vccd1 _3486_ sky130_fd_sc_hd__mux2_1
X_4454_ reg_data\[6\]\[2\] _1076_ _1048_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__and3_1
X_7173_ _3449_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__clkbuf_1
X_4385_ _1013_ vssd1 vssd1 vccd1 vccd1 rs2_mux\[3\] sky130_fd_sc_hd__clkinv_2
X_6124_ reg_data\[2\]\[27\] _2219_ _2396_ _2397_ reg_data\[11\]\[27\] vssd1 vssd1
+ vccd1 vccd1 _2697_ sky130_fd_sc_hd__a32o_1
X_6055_ reg_data\[25\]\[26\] _2370_ _2627_ _2628_ _2629_ vssd1 vssd1 vccd1 vccd1 _2630_
+ sky130_fd_sc_hd__a2111o_1
X_5006_ reg_data\[1\]\[9\] _1022_ _1109_ _1111_ reg_data\[15\]\[9\] vssd1 vssd1 vccd1
+ vccd1 _1615_ sky130_fd_sc_hd__a32o_1
X_9814_ clknet_leaf_39_i_clk rdata1\[30\] vssd1 vssd1 vccd1 vccd1 r_data1\[30\] sky130_fd_sc_hd__dfxtp_1
X_9745_ clknet_leaf_17_i_clk _0889_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6957_ _3248_ reg_data\[10\]\[22\] _3331_ vssd1 vssd1 vccd1 vccd1 _3334_ sky130_fd_sc_hd__mux2_1
X_5908_ reg_data\[22\]\[23\] _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__and3_1
X_9676_ clknet_leaf_29_i_clk _0820_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6888_ _3296_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__clkbuf_1
X_8627_ _4215_ vssd1 vssd1 vccd1 vccd1 _4238_ sky130_fd_sc_hd__buf_4
X_5839_ _1157_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__clkbuf_4
X_8558_ _4201_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__clkbuf_1
X_7509_ _3250_ reg_data\[21\]\[23\] _3625_ vssd1 vssd1 vccd1 vccd1 _3629_ sky130_fd_sc_hd__mux2_1
X_8489_ _3898_ reg_data\[18\]\[19\] _4155_ vssd1 vssd1 vccd1 vccd1 _4165_ sky130_fd_sc_hd__mux2_1
X_7860_ _3815_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__clkbuf_1
X_6811_ _3250_ reg_data\[22\]\[23\] _3244_ vssd1 vssd1 vccd1 vccd1 _3251_ sky130_fd_sc_hd__mux2_1
X_7791_ _3258_ reg_data\[26\]\[27\] _3771_ vssd1 vssd1 vccd1 vccd1 _3779_ sky130_fd_sc_hd__mux2_1
X_9530_ clknet_leaf_11_i_clk _0674_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6742_ i_data[1] vssd1 vssd1 vccd1 vccd1 _3204_ sky130_fd_sc_hd__clkbuf_4
X_9461_ clknet_leaf_32_i_clk _0605_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6673_ _3155_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__clkbuf_1
X_9392_ clknet_leaf_33_i_clk _0536_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_5624_ reg_data\[12\]\[19\] _1986_ _1606_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__and3_1
X_8412_ _4124_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__clkbuf_1
X_8343_ _3888_ reg_data\[16\]\[14\] _4083_ vssd1 vssd1 vccd1 vccd1 _4088_ sky130_fd_sc_hd__mux2_1
X_5555_ reg_data\[17\]\[18\] _2086_ _1108_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__and3_1
X_4506_ _1062_ _1128_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__and2_4
X_8274_ _3888_ reg_data\[15\]\[14\] _4046_ vssd1 vssd1 vccd1 vccd1 _4051_ sky130_fd_sc_hd__mux2_1
X_5486_ reg_data\[8\]\[16\] _1841_ _1842_ reg_data\[10\]\[16\] _2079_ vssd1 vssd1
+ vccd1 vccd1 _2080_ sky130_fd_sc_hd__a221o_1
X_4437_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__buf_4
X_7225_ reg_data\[6\]\[19\] _3168_ _3467_ vssd1 vssd1 vccd1 vccd1 _3477_ sky130_fd_sc_hd__mux2_1
X_7156_ _3440_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__clkbuf_1
X_6107_ reg_data\[17\]\[27\] _2372_ _1040_ vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__and3_1
X_4368_ _0999_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__clkbuf_4
X_7087_ _3403_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__clkbuf_1
X_6038_ reg_data\[14\]\[25\] _2301_ _1344_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__and3_1
X_7989_ i_data[16] vssd1 vssd1 vccd1 vccd1 _3892_ sky130_fd_sc_hd__clkbuf_4
X_9728_ clknet_leaf_5_i_clk _0872_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_9659_ clknet_leaf_4_i_clk _0803_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5340_ reg_data\[26\]\[14\] _1805_ _1806_ reg_data\[29\]\[14\] vssd1 vssd1 vccd1
+ vccd1 _1939_ sky130_fd_sc_hd__a22o_1
X_5271_ _1857_ _1861_ _1866_ _1871_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__or4_1
X_7010_ reg_data\[0\]\[15\] _3160_ _3356_ vssd1 vssd1 vccd1 vccd1 _3362_ sky130_fd_sc_hd__mux2_1
X_8961_ clknet_leaf_1_i_clk _0105_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_7912_ _3843_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__clkbuf_1
X_8892_ clknet_leaf_7_i_clk _0036_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_7843_ _3806_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__clkbuf_1
X_7774_ _3241_ reg_data\[26\]\[19\] _3760_ vssd1 vssd1 vccd1 vccd1 _3770_ sky130_fd_sc_hd__mux2_1
X_4986_ reg_data\[18\]\[9\] _1055_ _1483_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__and3_1
X_6725_ _3190_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__clkbuf_1
X_9513_ clknet_leaf_26_i_clk _0657_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_9444_ clknet_leaf_62_i_clk _0588_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_6656_ reg_data\[4\]\[7\] _3143_ _3129_ vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__mux2_1
X_6587_ _3099_ vssd1 vssd1 vccd1 vccd1 o_data2[14] sky130_fd_sc_hd__buf_2
X_9375_ clknet_leaf_1_i_clk _0519_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5607_ _2188_ _2192_ _2194_ _2196_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__or4_1
X_8326_ _3871_ reg_data\[16\]\[6\] _4072_ vssd1 vssd1 vccd1 vccd1 _4079_ sky130_fd_sc_hd__mux2_1
X_5538_ reg_data\[14\]\[17\] _1693_ _1958_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__and3_1
X_8257_ _3871_ reg_data\[15\]\[6\] _4035_ vssd1 vssd1 vccd1 vccd1 _4042_ sky130_fd_sc_hd__mux2_1
X_7208_ _3468_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
X_5469_ reg_data\[3\]\[16\] _1815_ _2060_ _2061_ _2062_ vssd1 vssd1 vccd1 vccd1 _2063_
+ sky130_fd_sc_hd__a2111o_1
X_8188_ _4005_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__clkbuf_1
X_7139_ reg_data\[7\]\[10\] _3149_ _3431_ vssd1 vssd1 vccd1 vccd1 _3432_ sky130_fd_sc_hd__mux2_1
X_4840_ reg_data\[25\]\[6\] _1141_ _1451_ _1452_ _1453_ vssd1 vssd1 vccd1 vccd1 _1454_
+ sky130_fd_sc_hd__a2111o_1
X_6510_ _3058_ vssd1 vssd1 vccd1 vccd1 o_data1[10] sky130_fd_sc_hd__buf_2
X_4771_ reg_data\[1\]\[5\] _1022_ _1109_ _1111_ reg_data\[15\]\[5\] vssd1 vssd1 vccd1
+ vccd1 _1388_ sky130_fd_sc_hd__a32o_1
X_7490_ _3231_ reg_data\[21\]\[14\] _3614_ vssd1 vssd1 vccd1 vccd1 _3619_ sky130_fd_sc_hd__mux2_1
X_6441_ reg_data\[5\]\[1\] _1085_ _2530_ vssd1 vssd1 vccd1 vccd1 _3002_ sky130_fd_sc_hd__and3_1
X_6372_ reg_data\[8\]\[31\] _2447_ _2448_ reg_data\[10\]\[31\] _2935_ vssd1 vssd1
+ vccd1 vccd1 _2936_ sky130_fd_sc_hd__a221o_1
X_9160_ clknet_leaf_46_i_clk _0304_ vssd1 vssd1 vccd1 vccd1 reg_data\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_8111_ _3861_ reg_data\[13\]\[1\] _3963_ vssd1 vssd1 vccd1 vccd1 _3965_ sky130_fd_sc_hd__mux2_1
X_5323_ reg_data\[3\]\[14\] _1770_ _1917_ _1920_ _1921_ vssd1 vssd1 vccd1 vccd1 _1922_
+ sky130_fd_sc_hd__a2111o_1
X_9091_ clknet_leaf_64_i_clk _0235_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8042_ _3861_ reg_data\[30\]\[1\] _3926_ vssd1 vssd1 vccd1 vccd1 _3928_ sky130_fd_sc_hd__mux2_1
X_5254_ reg_data\[21\]\[13\] _1766_ _1044_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__and3_1
X_5185_ _1100_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__clkbuf_4
X_8944_ clknet_leaf_37_i_clk _0088_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_8875_ clknet_leaf_43_i_clk _0019_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_7826_ _3225_ reg_data\[27\]\[11\] _3796_ vssd1 vssd1 vccd1 vccd1 _3798_ sky130_fd_sc_hd__mux2_1
X_7757_ _3761_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__clkbuf_1
X_4969_ reg_data\[12\]\[8\] _1354_ _1226_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__and3_1
X_6708_ i_data[24] vssd1 vssd1 vccd1 vccd1 _3179_ sky130_fd_sc_hd__clkbuf_4
X_7688_ _3222_ reg_data\[25\]\[10\] _3724_ vssd1 vssd1 vccd1 vccd1 _3725_ sky130_fd_sc_hd__mux2_1
X_9427_ clknet_leaf_35_i_clk _0571_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6639_ _3132_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__clkbuf_1
X_9358_ clknet_leaf_39_i_clk _0502_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_8309_ _3923_ reg_data\[15\]\[31\] _4034_ vssd1 vssd1 vccd1 vccd1 _4069_ sky130_fd_sc_hd__mux2_1
X_9289_ clknet_leaf_58_i_clk _0433_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_44_i_clk clknet_3_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_6990_ _3351_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__clkbuf_1
X_5941_ reg_data\[17\]\[24\] _2372_ _1708_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__and3_1
X_5872_ _1227_ vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_59_i_clk clknet_3_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_8660_ reg_data\[19\]\[3\] _3135_ _4252_ vssd1 vssd1 vccd1 vccd1 _4256_ sky130_fd_sc_hd__mux2_1
X_8591_ _4219_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__clkbuf_1
X_7611_ _3214_ reg_data\[24\]\[6\] _3677_ vssd1 vssd1 vccd1 vccd1 _3684_ sky130_fd_sc_hd__mux2_1
X_4823_ reg_data\[12\]\[6\] _1381_ _1128_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__and3_1
X_7542_ reg_data\[23\]\[6\] _3141_ _3640_ vssd1 vssd1 vccd1 vccd1 _3647_ sky130_fd_sc_hd__mux2_1
X_4754_ reg_data\[18\]\[5\] _1055_ _1064_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__and3_1
X_7473_ _3214_ reg_data\[21\]\[6\] _3603_ vssd1 vssd1 vccd1 vccd1 _3610_ sky130_fd_sc_hd__mux2_1
X_4685_ reg_data\[24\]\[3\] _1225_ _1228_ reg_data\[28\]\[3\] _1304_ vssd1 vssd1 vccd1
+ vccd1 _1305_ sky130_fd_sc_hd__a221o_1
X_9212_ clknet_leaf_7_i_clk _0356_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6424_ reg_data\[27\]\[0\] _1198_ _2983_ _2984_ _2985_ vssd1 vssd1 vccd1 vccd1 _2986_
+ sky130_fd_sc_hd__a2111o_1
X_9143_ clknet_leaf_14_i_clk _0287_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6355_ reg_data\[30\]\[31\] _1146_ _1163_ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__and3_1
X_9074_ clknet_leaf_17_i_clk _0218_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6286_ reg_data\[2\]\[30\] _1021_ _2396_ _2397_ reg_data\[11\]\[30\] vssd1 vssd1
+ vccd1 vccd1 _2853_ sky130_fd_sc_hd__a32o_1
X_5306_ reg_data\[1\]\[13\] _1904_ _1905_ reg_data\[15\]\[13\] vssd1 vssd1 vccd1 vccd1
+ _1906_ sky130_fd_sc_hd__a22o_1
X_8025_ _3916_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__clkbuf_1
X_5237_ reg_data\[1\]\[12\] _1298_ _1299_ reg_data\[15\]\[12\] vssd1 vssd1 vccd1 vccd1
+ _1839_ sky130_fd_sc_hd__a22o_1
X_5168_ reg_data\[18\]\[12\] _1656_ _1483_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__and3_1
X_5099_ reg_data\[24\]\[10\] _1225_ _1228_ reg_data\[28\]\[10\] _1704_ vssd1 vssd1
+ vccd1 vccd1 _1705_ sky130_fd_sc_hd__a221o_1
X_8927_ clknet_leaf_77_i_clk _0071_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8858_ clknet_leaf_12_i_clk _0002_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_7809_ _3208_ reg_data\[27\]\[3\] _3785_ vssd1 vssd1 vccd1 vccd1 _3789_ sky130_fd_sc_hd__mux2_1
X_8789_ _4323_ vssd1 vssd1 vccd1 vccd1 _4324_ sky130_fd_sc_hd__buf_4
X_4470_ _1050_ _1066_ _1078_ _1092_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__or4_2
X_6140_ reg_data\[3\]\[27\] _2421_ _2709_ _2710_ _2711_ vssd1 vssd1 vccd1 vccd1 _2712_
+ sky130_fd_sc_hd__a2111o_1
X_6071_ reg_data\[1\]\[26\] _2336_ _2399_ _2400_ reg_data\[15\]\[26\] vssd1 vssd1
+ vccd1 vccd1 _2646_ sky130_fd_sc_hd__a32o_1
X_5022_ reg_data\[20\]\[9\] _1629_ _1180_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__and3_1
X_9830_ clknet_leaf_50_i_clk rdata2\[14\] vssd1 vssd1 vccd1 vccd1 r_data2\[14\] sky130_fd_sc_hd__dfxtp_1
X_6973_ _3264_ reg_data\[10\]\[30\] _3308_ vssd1 vssd1 vccd1 vccd1 _3342_ sky130_fd_sc_hd__mux2_1
X_9761_ clknet_leaf_1_i_clk _0905_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5924_ reg_data\[7\]\[23\] _2433_ _2501_ _2502_ _2503_ vssd1 vssd1 vccd1 vccd1 _2504_
+ sky130_fd_sc_hd__a2111o_1
X_8712_ reg_data\[19\]\[28\] _3187_ _4274_ vssd1 vssd1 vccd1 vccd1 _4283_ sky130_fd_sc_hd__mux2_1
X_9692_ clknet_leaf_76_i_clk _0836_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_8643_ _4246_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__clkbuf_1
X_5855_ reg_data\[7\]\[22\] _2433_ _2434_ _2435_ _2436_ vssd1 vssd1 vccd1 vccd1 _2437_
+ sky130_fd_sc_hd__a2111o_1
X_4806_ reg_data\[26\]\[5\] _1230_ _1232_ reg_data\[29\]\[5\] vssd1 vssd1 vccd1 vccd1
+ _1422_ sky130_fd_sc_hd__a22o_1
X_8574_ reg_data\[1\]\[27\] _3185_ _4202_ vssd1 vssd1 vccd1 vccd1 _4210_ sky130_fd_sc_hd__mux2_1
X_5786_ _2369_ vssd1 vssd1 vccd1 vccd1 rdata2\[21\] sky130_fd_sc_hd__clkbuf_1
X_7525_ _3266_ reg_data\[21\]\[31\] _3602_ vssd1 vssd1 vccd1 vccd1 _3637_ sky130_fd_sc_hd__mux2_1
X_4737_ reg_data\[12\]\[4\] _1354_ _1226_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__and3_1
X_7456_ _3599_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__clkbuf_1
X_4668_ reg_data\[14\]\[3\] _1186_ _1164_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__and3_1
X_6407_ reg_data\[25\]\[0\] _2416_ _2966_ _2967_ _2968_ vssd1 vssd1 vccd1 vccd1 _2969_
+ sky130_fd_sc_hd__a2111o_1
X_7387_ reg_data\[3\]\[31\] _3193_ _3528_ vssd1 vssd1 vccd1 vccd1 _3563_ sky130_fd_sc_hd__mux2_1
X_4599_ _1220_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__clkbuf_4
X_9126_ clknet_leaf_47_i_clk _0270_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6338_ _2890_ _2894_ _2898_ _2902_ vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__or4_2
X_6269_ reg_data\[17\]\[30\] _2372_ _1040_ vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__and3_1
X_9057_ clknet_leaf_5_i_clk _0201_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_8008_ i_data[22] vssd1 vssd1 vccd1 vccd1 _3905_ sky130_fd_sc_hd__clkbuf_4
X_5640_ reg_data\[22\]\[19\] _1679_ _1622_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__and3_1
X_5571_ reg_data\[23\]\[18\] _1787_ _1788_ reg_data\[19\]\[18\] vssd1 vssd1 vccd1
+ vccd1 _2162_ sky130_fd_sc_hd__a22o_1
X_7310_ _3522_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__clkbuf_1
X_4522_ rs2_mux\[0\] _1006_ rs2_mux\[2\] _1013_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__and4_4
X_8290_ _4059_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__clkbuf_1
X_7241_ _3485_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__clkbuf_1
X_4453_ _1067_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__buf_2
X_7172_ reg_data\[7\]\[26\] _3183_ _3442_ vssd1 vssd1 vccd1 vccd1 _3449_ sky130_fd_sc_hd__mux2_1
X_4384_ _0994_ _0996_ _1011_ _1012_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__a31o_2
X_6123_ reg_data\[23\]\[27\] _2393_ _2394_ reg_data\[19\]\[27\] vssd1 vssd1 vccd1
+ vccd1 _2696_ sky130_fd_sc_hd__a22o_1
X_6054_ reg_data\[17\]\[26\] _2086_ _1238_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__and3_1
X_5005_ reg_data\[2\]\[9\] _1613_ _1104_ _1106_ reg_data\[11\]\[9\] vssd1 vssd1 vccd1
+ vccd1 _1614_ sky130_fd_sc_hd__a32o_1
X_9813_ clknet_leaf_36_i_clk rdata1\[29\] vssd1 vssd1 vccd1 vccd1 r_data1\[29\] sky130_fd_sc_hd__dfxtp_1
X_9744_ clknet_leaf_19_i_clk _0888_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6956_ _3333_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__clkbuf_1
X_5907_ _2487_ vssd1 vssd1 vccd1 vccd1 rdata1\[23\] sky130_fd_sc_hd__clkbuf_1
X_6887_ reg_data\[2\]\[22\] _3175_ _3293_ vssd1 vssd1 vccd1 vccd1 _3296_ sky130_fd_sc_hd__mux2_1
X_9675_ clknet_leaf_44_i_clk _0819_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5838_ reg_data\[25\]\[22\] _2416_ _2417_ _2418_ _2419_ vssd1 vssd1 vccd1 vccd1 _2420_
+ sky130_fd_sc_hd__a2111o_1
X_8626_ _4237_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__clkbuf_1
X_5769_ reg_data\[4\]\[21\] _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__and3_1
X_8557_ reg_data\[1\]\[19\] _3168_ _4191_ vssd1 vssd1 vccd1 vccd1 _4201_ sky130_fd_sc_hd__mux2_1
X_7508_ _3628_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__clkbuf_1
X_8488_ _4164_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__clkbuf_1
X_7439_ _3250_ reg_data\[20\]\[23\] _3587_ vssd1 vssd1 vccd1 vccd1 _3591_ sky130_fd_sc_hd__mux2_1
X_9109_ clknet_leaf_16_i_clk _0253_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6810_ i_data[23] vssd1 vssd1 vccd1 vccd1 _3250_ sky130_fd_sc_hd__buf_2
X_7790_ _3778_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__clkbuf_1
X_6741_ _3203_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__clkbuf_1
X_9460_ clknet_leaf_32_i_clk _0604_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6672_ reg_data\[4\]\[12\] _3154_ _3150_ vssd1 vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__mux2_1
X_9391_ clknet_leaf_32_i_clk _0535_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_5623_ reg_data\[14\]\[19\] _1867_ _2156_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__and3_1
X_8411_ _3888_ reg_data\[17\]\[14\] _4119_ vssd1 vssd1 vccd1 vccd1 _4124_ sky130_fd_sc_hd__mux2_1
X_8342_ _4087_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__clkbuf_1
X_5554_ reg_data\[21\]\[18\] _1766_ _1044_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__and3_1
X_4505_ _1083_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__clkbuf_4
X_8273_ _4050_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__clkbuf_1
X_5485_ reg_data\[16\]\[16\] _1843_ _1844_ reg_data\[9\]\[16\] vssd1 vssd1 vccd1 vccd1
+ _2079_ sky130_fd_sc_hd__a22o_1
X_4436_ _1015_ _1026_ rs1_mux\[2\] _1033_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__and4_4
X_7224_ _3476_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
X_4367_ _0995_ i_rs2[4] _0996_ _0998_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__o31a_2
X_7155_ reg_data\[7\]\[18\] _3166_ _3431_ vssd1 vssd1 vccd1 vccd1 _3440_ sky130_fd_sc_hd__mux2_1
X_6106_ reg_data\[22\]\[27\] _2143_ _2256_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__and3_1
X_7086_ _3239_ reg_data\[8\]\[18\] _3394_ vssd1 vssd1 vccd1 vccd1 _3403_ sky130_fd_sc_hd__mux2_1
X_6037_ reg_data\[13\]\[25\] _2183_ _2299_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__and3_1
X_7988_ _3891_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__clkbuf_1
X_6939_ _3324_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__clkbuf_1
X_9727_ clknet_leaf_4_i_clk _0871_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_9658_ clknet_leaf_11_i_clk _0802_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8609_ _3882_ reg_data\[12\]\[11\] _4227_ vssd1 vssd1 vccd1 vccd1 _4229_ sky130_fd_sc_hd__mux2_1
X_9589_ clknet_leaf_37_i_clk _0733_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_5270_ reg_data\[7\]\[13\] _1780_ _1868_ _1869_ _1870_ vssd1 vssd1 vccd1 vccd1 _1871_
+ sky130_fd_sc_hd__a2111o_1
X_8960_ clknet_leaf_74_i_clk _0104_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7911_ _3241_ reg_data\[28\]\[19\] _3833_ vssd1 vssd1 vccd1 vccd1 _3843_ sky130_fd_sc_hd__mux2_1
X_8891_ clknet_leaf_2_i_clk _0035_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_7842_ _3241_ reg_data\[27\]\[19\] _3796_ vssd1 vssd1 vccd1 vccd1 _3806_ sky130_fd_sc_hd__mux2_1
X_7773_ _3769_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__clkbuf_1
X_4985_ reg_data\[25\]\[9\] _1037_ _1591_ _1592_ _1593_ vssd1 vssd1 vccd1 vccd1 _1594_
+ sky130_fd_sc_hd__a2111o_1
X_6724_ reg_data\[4\]\[29\] _3189_ _3171_ vssd1 vssd1 vccd1 vccd1 _3190_ sky130_fd_sc_hd__mux2_1
X_9512_ clknet_leaf_45_i_clk _0656_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_9443_ clknet_leaf_62_i_clk _0587_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_0__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_6655_ i_data[7] vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__buf_2
X_9374_ clknet_leaf_77_i_clk _0518_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_5606_ reg_data\[24\]\[18\] _1847_ _1848_ reg_data\[28\]\[18\] _2195_ vssd1 vssd1
+ vccd1 vccd1 _2196_ sky130_fd_sc_hd__a221o_1
X_6586_ r_data2\[14\] _3094_ vssd1 vssd1 vccd1 vccd1 _3099_ sky130_fd_sc_hd__and2_1
X_5537_ reg_data\[13\]\[17\] _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__and3_1
X_8325_ _4078_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__clkbuf_1
X_8256_ _4041_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__clkbuf_1
X_7207_ reg_data\[6\]\[10\] _3149_ _3467_ vssd1 vssd1 vccd1 vccd1 _3468_ sky130_fd_sc_hd__mux2_1
X_5468_ reg_data\[20\]\[16\] _1629_ _1743_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__and3_1
X_5399_ reg_data\[8\]\[15\] _1797_ _1798_ reg_data\[10\]\[15\] _1995_ vssd1 vssd1
+ vccd1 vccd1 _1996_ sky130_fd_sc_hd__a221o_1
X_8187_ _3869_ reg_data\[14\]\[5\] _3999_ vssd1 vssd1 vccd1 vccd1 _4005_ sky130_fd_sc_hd__mux2_1
X_4419_ _1038_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__buf_2
X_7138_ _3419_ vssd1 vssd1 vccd1 vccd1 _3431_ sky130_fd_sc_hd__buf_4
X_7069_ _3382_ vssd1 vssd1 vccd1 vccd1 _3394_ sky130_fd_sc_hd__buf_4
X_4770_ reg_data\[2\]\[5\] _1103_ _1104_ _1106_ reg_data\[11\]\[5\] vssd1 vssd1 vccd1
+ vccd1 _1387_ sky130_fd_sc_hd__a32o_1
X_6440_ reg_data\[4\]\[1\] _1072_ _1060_ vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__and3_1
X_6371_ reg_data\[16\]\[31\] _2449_ _2450_ reg_data\[9\]\[31\] vssd1 vssd1 vccd1 vccd1
+ _2935_ sky130_fd_sc_hd__a22o_1
X_8110_ _3964_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__clkbuf_1
X_5322_ reg_data\[20\]\[14\] _1597_ _1315_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__and3_1
X_9090_ clknet_leaf_66_i_clk _0234_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8041_ _3927_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__clkbuf_1
X_5253_ reg_data\[22\]\[13\] _1536_ _1651_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__and3_1
X_5184_ _1098_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__buf_4
X_8943_ clknet_leaf_37_i_clk _0087_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_8874_ clknet_leaf_41_i_clk _0018_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_7825_ _3797_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__clkbuf_1
X_7756_ _3222_ reg_data\[26\]\[10\] _3760_ vssd1 vssd1 vccd1 vccd1 _3761_ sky130_fd_sc_hd__mux2_1
X_4968_ reg_data\[14\]\[8\] _1189_ _1193_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__and3_1
X_6707_ _3178_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__clkbuf_1
X_7687_ _3712_ vssd1 vssd1 vccd1 vccd1 _3724_ sky130_fd_sc_hd__buf_4
X_4899_ reg_data\[21\]\[7\] _1509_ _1510_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__and3_1
X_9426_ clknet_leaf_34_i_clk _0570_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6638_ reg_data\[4\]\[1\] _3131_ _3129_ vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__mux2_1
X_9357_ clknet_leaf_50_i_clk _0501_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_8308_ _4068_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__clkbuf_1
X_6569_ r_data2\[6\] _3083_ vssd1 vssd1 vccd1 vccd1 _3090_ sky130_fd_sc_hd__and2_1
X_9288_ clknet_leaf_53_i_clk _0432_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_8239_ _3921_ reg_data\[14\]\[30\] _3998_ vssd1 vssd1 vccd1 vccd1 _4032_ sky130_fd_sc_hd__mux2_1
X_5940_ reg_data\[22\]\[24\] _2143_ _2256_ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__and3_1
X_5871_ _1224_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__clkbuf_4
X_7610_ _3683_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__clkbuf_1
X_8590_ _3863_ reg_data\[12\]\[2\] _4216_ vssd1 vssd1 vccd1 vccd1 _4219_ sky130_fd_sc_hd__mux2_1
X_4822_ reg_data\[14\]\[6\] _1253_ _1379_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__and3_1
X_7541_ _3646_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__clkbuf_1
X_4753_ reg_data\[25\]\[5\] _1037_ _1367_ _1368_ _1369_ vssd1 vssd1 vccd1 vccd1 _1370_
+ sky130_fd_sc_hd__a2111o_1
X_7472_ _3609_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__clkbuf_1
X_4684_ reg_data\[26\]\[3\] _1230_ _1232_ reg_data\[29\]\[3\] vssd1 vssd1 vccd1 vccd1
+ _1304_ sky130_fd_sc_hd__a22o_1
X_6423_ reg_data\[1\]\[0\] _2510_ _2511_ reg_data\[15\]\[0\] vssd1 vssd1 vccd1 vccd1
+ _2985_ sky130_fd_sc_hd__a22o_1
X_9211_ clknet_leaf_6_i_clk _0355_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_9142_ clknet_leaf_14_i_clk _0286_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6354_ reg_data\[18\]\[31\] _2422_ _1167_ vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__and3_1
X_9073_ clknet_leaf_18_i_clk _0217_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6285_ reg_data\[23\]\[30\] _2393_ _2394_ reg_data\[19\]\[30\] vssd1 vssd1 vccd1
+ vccd1 _2852_ sky130_fd_sc_hd__a22o_1
X_5305_ _1203_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__buf_4
X_8024_ _3915_ reg_data\[9\]\[27\] _3901_ vssd1 vssd1 vccd1 vccd1 _3916_ sky130_fd_sc_hd__mux2_1
X_5236_ reg_data\[2\]\[12\] _1837_ _1295_ _1296_ reg_data\[11\]\[12\] vssd1 vssd1
+ vccd1 vccd1 _1838_ sky130_fd_sc_hd__a32o_1
X_5167_ _1053_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__buf_4
X_5098_ reg_data\[26\]\[10\] _1230_ _1232_ reg_data\[29\]\[10\] vssd1 vssd1 vccd1
+ vccd1 _1704_ sky130_fd_sc_hd__a22o_1
X_8926_ clknet_leaf_76_i_clk _0070_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8857_ clknet_leaf_11_i_clk _0001_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8788_ _3307_ _3638_ vssd1 vssd1 vccd1 vccd1 _4323_ sky130_fd_sc_hd__and2_4
X_7808_ _3788_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__clkbuf_1
X_7739_ _3206_ reg_data\[26\]\[2\] _3749_ vssd1 vssd1 vccd1 vccd1 _3752_ sky130_fd_sc_hd__mux2_1
X_9409_ clknet_leaf_72_i_clk _0553_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6070_ reg_data\[2\]\[26\] _2219_ _2396_ _2397_ reg_data\[11\]\[26\] vssd1 vssd1
+ vccd1 vccd1 _2645_ sky130_fd_sc_hd__a32o_1
X_5021_ _1138_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__buf_2
X_9760_ clknet_leaf_76_i_clk _0904_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8711_ _4282_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__clkbuf_1
X_6972_ _3341_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__clkbuf_1
X_5923_ reg_data\[12\]\[23\] _1960_ _2016_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__and3_1
X_9691_ clknet_leaf_76_i_clk _0835_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_8642_ _3915_ reg_data\[12\]\[27\] _4238_ vssd1 vssd1 vccd1 vccd1 _4246_ sky130_fd_sc_hd__mux2_1
X_5854_ reg_data\[12\]\[22\] _1960_ _2016_ vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__and3_1
X_8573_ _4209_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__clkbuf_1
X_4805_ reg_data\[8\]\[5\] _1214_ _1217_ reg_data\[10\]\[5\] _1420_ vssd1 vssd1 vccd1
+ vccd1 _1421_ sky130_fd_sc_hd__a221o_1
X_7524_ _3636_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__clkbuf_1
X_5785_ _2360_ _2364_ _2366_ _2368_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__or4_1
X_4736_ _1000_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__buf_2
X_7455_ _3266_ reg_data\[20\]\[31\] _3564_ vssd1 vssd1 vccd1 vccd1 _3599_ sky130_fd_sc_hd__mux2_1
X_4667_ reg_data\[0\]\[3\] _1174_ _1282_ _1284_ _1286_ vssd1 vssd1 vccd1 vccd1 _1287_
+ sky130_fd_sc_hd__a2111o_1
X_7386_ _3562_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__clkbuf_1
X_6406_ reg_data\[21\]\[0\] _1162_ _1510_ vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__and3_1
X_6337_ reg_data\[7\]\[31\] _2386_ _2899_ _2900_ _2901_ vssd1 vssd1 vccd1 vccd1 _2902_
+ sky130_fd_sc_hd__a2111o_1
X_4598_ _1000_ _1139_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__and2_4
X_9125_ clknet_leaf_63_i_clk _0269_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6268_ reg_data\[22\]\[30\] _1097_ _1047_ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__and3_1
X_9056_ clknet_leaf_5_i_clk _0200_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6199_ reg_data\[13\]\[28\] _1177_ _2299_ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__and3_1
X_5219_ _1173_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__clkbuf_4
X_8007_ _3904_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__clkbuf_1
X_8909_ clknet_leaf_28_i_clk _0053_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_9889_ clknet_leaf_38_i_clk _0959_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_43_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_58_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5570_ _2147_ _2151_ _2155_ _2160_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__or4_2
X_4521_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__buf_2
X_7240_ reg_data\[6\]\[26\] _3183_ _3478_ vssd1 vssd1 vccd1 vccd1 _3485_ sky130_fd_sc_hd__mux2_1
X_4452_ reg_data\[5\]\[2\] _1074_ _1044_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__and3_1
X_7171_ _3448_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__clkbuf_1
X_4383_ _0994_ rs2\[3\] vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__nor2_1
X_6122_ _2682_ _2686_ _2690_ _2694_ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__or4_4
X_6053_ reg_data\[21\]\[26\] _2372_ _1043_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__and3_1
X_5004_ _1089_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__buf_4
X_9812_ clknet_leaf_32_i_clk rdata1\[28\] vssd1 vssd1 vccd1 vccd1 r_data1\[28\] sky130_fd_sc_hd__dfxtp_1
X_9743_ clknet_leaf_23_i_clk _0887_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6955_ _3246_ reg_data\[10\]\[21\] _3331_ vssd1 vssd1 vccd1 vccd1 _3333_ sky130_fd_sc_hd__mux2_1
X_5906_ _2478_ _2482_ _2484_ _2486_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__or4_1
X_9674_ clknet_leaf_43_i_clk _0818_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8625_ _3898_ reg_data\[12\]\[19\] _4227_ vssd1 vssd1 vccd1 vccd1 _4237_ sky130_fd_sc_hd__mux2_1
X_6886_ _3295_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__clkbuf_1
X_5837_ reg_data\[17\]\[22\] _2117_ _1148_ vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__and3_1
X_5768_ reg_data\[6\]\[21\] _1951_ _2237_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__and3_1
X_8556_ _4200_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__clkbuf_1
X_7507_ _3248_ reg_data\[21\]\[22\] _3625_ vssd1 vssd1 vccd1 vccd1 _3628_ sky130_fd_sc_hd__mux2_1
X_8487_ _3896_ reg_data\[18\]\[18\] _4155_ vssd1 vssd1 vccd1 vccd1 _4164_ sky130_fd_sc_hd__mux2_1
X_4719_ reg_data\[17\]\[4\] _1272_ _1148_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__and3_1
X_7438_ _3590_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__clkbuf_1
X_5699_ _0997_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__buf_2
X_7369_ reg_data\[3\]\[22\] _3175_ _3551_ vssd1 vssd1 vccd1 vccd1 _3554_ sky130_fd_sc_hd__mux2_1
X_9108_ clknet_leaf_18_i_clk _0252_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_9039_ clknet_leaf_32_i_clk _0183_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6740_ _3195_ reg_data\[22\]\[0\] _3202_ vssd1 vssd1 vccd1 vccd1 _3203_ sky130_fd_sc_hd__mux2_1
X_6671_ i_data[12] vssd1 vssd1 vccd1 vccd1 _3154_ sky130_fd_sc_hd__buf_2
X_9390_ clknet_leaf_39_i_clk _0534_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_5622_ reg_data\[0\]\[19\] _1775_ _2208_ _2209_ _2210_ vssd1 vssd1 vccd1 vccd1 _2211_
+ sky130_fd_sc_hd__a2111o_1
X_8410_ _4123_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__clkbuf_1
X_5553_ reg_data\[22\]\[18\] _2143_ _1651_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__and3_1
X_8341_ _3886_ reg_data\[16\]\[13\] _4083_ vssd1 vssd1 vccd1 vccd1 _4087_ sky130_fd_sc_hd__mux2_1
X_4504_ _1126_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__clkbuf_4
X_8272_ _3886_ reg_data\[15\]\[13\] _4046_ vssd1 vssd1 vccd1 vccd1 _4050_ sky130_fd_sc_hd__mux2_1
X_5484_ reg_data\[27\]\[16\] _1833_ _2075_ _2076_ _2077_ vssd1 vssd1 vccd1 vccd1 _2078_
+ sky130_fd_sc_hd__a2111o_1
X_7223_ reg_data\[6\]\[18\] _3166_ _3467_ vssd1 vssd1 vccd1 vccd1 _3476_ sky130_fd_sc_hd__mux2_1
X_4435_ _1034_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__clkbuf_4
X_4366_ _0995_ _0996_ _0997_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__o21ai_1
X_7154_ _3439_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__clkbuf_1
X_6105_ _2678_ vssd1 vssd1 vccd1 vccd1 rdata2\[26\] sky130_fd_sc_hd__clkbuf_1
X_7085_ _3402_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__clkbuf_1
X_6036_ reg_data\[0\]\[25\] _2427_ _2609_ _2610_ _2611_ vssd1 vssd1 vccd1 vccd1 _2612_
+ sky130_fd_sc_hd__a2111o_1
X_7987_ _3890_ reg_data\[9\]\[15\] _3880_ vssd1 vssd1 vccd1 vccd1 _3891_ sky130_fd_sc_hd__mux2_1
X_6938_ _3229_ reg_data\[10\]\[13\] _3320_ vssd1 vssd1 vccd1 vccd1 _3324_ sky130_fd_sc_hd__mux2_1
X_9726_ clknet_leaf_4_i_clk _0870_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_9657_ clknet_leaf_12_i_clk _0801_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6869_ _3286_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__clkbuf_1
X_9588_ clknet_leaf_32_i_clk _0732_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_8608_ _4228_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__clkbuf_1
X_8539_ reg_data\[1\]\[10\] _3149_ _4191_ vssd1 vssd1 vccd1 vccd1 _4192_ sky130_fd_sc_hd__mux2_1
X_7910_ _3842_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__clkbuf_1
X_8890_ clknet_leaf_9_i_clk _0034_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_7841_ _3805_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__clkbuf_1
X_7772_ _3239_ reg_data\[26\]\[18\] _3760_ vssd1 vssd1 vccd1 vccd1 _3769_ sky130_fd_sc_hd__mux2_1
X_4984_ reg_data\[21\]\[9\] _1480_ _1240_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__and3_1
X_6723_ i_data[29] vssd1 vssd1 vccd1 vccd1 _3189_ sky130_fd_sc_hd__buf_4
X_9511_ clknet_leaf_8_i_clk _0655_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_9442_ clknet_leaf_62_i_clk _0586_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6654_ _3142_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__clkbuf_1
X_5605_ reg_data\[26\]\[18\] _1849_ _1850_ reg_data\[29\]\[18\] vssd1 vssd1 vccd1
+ vccd1 _2195_ sky130_fd_sc_hd__a22o_1
X_6585_ _3098_ vssd1 vssd1 vccd1 vccd1 o_data2[13] sky130_fd_sc_hd__buf_2
X_9373_ clknet_leaf_1_i_clk _0517_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_5536_ reg_data\[0\]\[17\] _1821_ _2125_ _2126_ _2127_ vssd1 vssd1 vccd1 vccd1 _2128_
+ sky130_fd_sc_hd__a2111o_1
X_8324_ _3869_ reg_data\[16\]\[5\] _4072_ vssd1 vssd1 vccd1 vccd1 _4078_ sky130_fd_sc_hd__mux2_1
X_8255_ _3869_ reg_data\[15\]\[5\] _4035_ vssd1 vssd1 vccd1 vccd1 _4041_ sky130_fd_sc_hd__mux2_1
X_5467_ reg_data\[30\]\[16\] _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__and3_1
X_7206_ _3455_ vssd1 vssd1 vccd1 vccd1 _3467_ sky130_fd_sc_hd__buf_6
X_4418_ reg_data\[17\]\[2\] _1039_ _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__and3_1
X_5398_ reg_data\[16\]\[15\] _1799_ _1800_ reg_data\[9\]\[15\] vssd1 vssd1 vccd1 vccd1
+ _1995_ sky130_fd_sc_hd__a22o_1
X_8186_ _4004_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__clkbuf_1
X_7137_ _3430_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
X_7068_ _3393_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
X_6019_ reg_data\[16\]\[25\] _2405_ _2406_ reg_data\[9\]\[25\] vssd1 vssd1 vccd1 vccd1
+ _2596_ sky130_fd_sc_hd__a22o_1
X_9709_ clknet_leaf_40_i_clk _0853_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6370_ reg_data\[27\]\[31\] _2439_ _2931_ _2932_ _2933_ vssd1 vssd1 vccd1 vccd1 _2934_
+ sky130_fd_sc_hd__a2111o_1
X_5321_ reg_data\[30\]\[14\] _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__and3_1
X_8040_ _3857_ reg_data\[30\]\[0\] _3926_ vssd1 vssd1 vccd1 vccd1 _3927_ sky130_fd_sc_hd__mux2_1
X_5252_ _1853_ vssd1 vssd1 vccd1 vccd1 rdata2\[12\] sky130_fd_sc_hd__clkbuf_1
X_5183_ _1095_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__buf_4
X_8942_ clknet_leaf_39_i_clk _0086_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_8873_ clknet_leaf_41_i_clk _0017_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_7824_ _3222_ reg_data\[27\]\[10\] _3796_ vssd1 vssd1 vccd1 vccd1 _3797_ sky130_fd_sc_hd__mux2_1
X_7755_ _3748_ vssd1 vssd1 vccd1 vccd1 _3760_ sky130_fd_sc_hd__buf_4
X_4967_ reg_data\[13\]\[8\] _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__and3_1
X_6706_ reg_data\[4\]\[23\] _3177_ _3171_ vssd1 vssd1 vccd1 vccd1 _3178_ sky130_fd_sc_hd__mux2_1
X_4898_ _1144_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__buf_4
X_7686_ _3723_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__clkbuf_1
X_9425_ clknet_leaf_35_i_clk _0569_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6637_ i_data[1] vssd1 vssd1 vccd1 vccd1 _3131_ sky130_fd_sc_hd__clkbuf_4
X_6568_ _3089_ vssd1 vssd1 vccd1 vccd1 o_data2[5] sky130_fd_sc_hd__buf_2
X_9356_ clknet_leaf_50_i_clk _0500_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8307_ _3921_ reg_data\[15\]\[30\] _4034_ vssd1 vssd1 vccd1 vccd1 _4068_ sky130_fd_sc_hd__mux2_1
X_5519_ reg_data\[26\]\[17\] _1805_ _1806_ reg_data\[29\]\[17\] vssd1 vssd1 vccd1
+ vccd1 _2112_ sky130_fd_sc_hd__a22o_1
X_6499_ _3052_ vssd1 vssd1 vccd1 vccd1 o_data1[5] sky130_fd_sc_hd__buf_2
X_9287_ clknet_leaf_52_i_clk _0431_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8238_ _4031_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__clkbuf_1
X_8169_ _3919_ reg_data\[13\]\[29\] _3985_ vssd1 vssd1 vccd1 vccd1 _3995_ sky130_fd_sc_hd__mux2_1
X_5870_ reg_data\[8\]\[22\] _2447_ _2448_ reg_data\[10\]\[22\] _2451_ vssd1 vssd1
+ vccd1 vccd1 _2452_ sky130_fd_sc_hd__a221o_1
X_4821_ reg_data\[0\]\[6\] _1070_ _1433_ _1434_ _1435_ vssd1 vssd1 vccd1 vccd1 _1436_
+ sky130_fd_sc_hd__a2111o_1
X_7540_ reg_data\[23\]\[5\] _3139_ _3640_ vssd1 vssd1 vccd1 vccd1 _3646_ sky130_fd_sc_hd__mux2_1
X_4752_ reg_data\[21\]\[5\] _1046_ _1240_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__and3_1
X_4683_ reg_data\[8\]\[3\] _1214_ _1217_ reg_data\[10\]\[3\] _1302_ vssd1 vssd1 vccd1
+ vccd1 _1303_ sky130_fd_sc_hd__a221o_1
X_7471_ _3212_ reg_data\[21\]\[5\] _3603_ vssd1 vssd1 vccd1 vccd1 _3609_ sky130_fd_sc_hd__mux2_1
X_6422_ reg_data\[2\]\[0\] _1001_ _2507_ _2508_ reg_data\[11\]\[0\] vssd1 vssd1 vccd1
+ vccd1 _2984_ sky130_fd_sc_hd__a32o_1
X_9210_ clknet_leaf_9_i_clk _0354_ vssd1 vssd1 vccd1 vccd1 reg_data\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_9141_ clknet_leaf_16_i_clk _0285_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6353_ _2913_ _2914_ _2915_ _2916_ vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__or4_1
X_9072_ clknet_leaf_19_i_clk _0216_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6284_ _2838_ _2842_ _2846_ _2850_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__or4_4
X_5304_ _1202_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__buf_4
X_8023_ i_data[27] vssd1 vssd1 vccd1 vccd1 _3915_ sky130_fd_sc_hd__clkbuf_4
X_5235_ _1001_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__clkbuf_4
X_5166_ reg_data\[25\]\[12\] _1764_ _1765_ _1767_ _1768_ vssd1 vssd1 vccd1 vccd1 _1769_
+ sky130_fd_sc_hd__a2111o_1
X_5097_ reg_data\[8\]\[10\] _1214_ _1217_ reg_data\[10\]\[10\] _1702_ vssd1 vssd1
+ vccd1 vccd1 _1703_ sky130_fd_sc_hd__a221o_1
X_8925_ clknet_leaf_0_i_clk _0069_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_8856_ clknet_leaf_14_i_clk _0000_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_5999_ reg_data\[17\]\[25\] _2372_ _1708_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__and3_1
X_8787_ _4322_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__clkbuf_1
X_7807_ _3206_ reg_data\[27\]\[2\] _3785_ vssd1 vssd1 vccd1 vccd1 _3788_ sky130_fd_sc_hd__mux2_1
X_7738_ _3751_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__clkbuf_1
X_7669_ _3204_ reg_data\[25\]\[1\] _3713_ vssd1 vssd1 vccd1 vccd1 _3715_ sky130_fd_sc_hd__mux2_1
X_9408_ clknet_leaf_70_i_clk _0552_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_9339_ clknet_leaf_71_i_clk _0483_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5020_ reg_data\[30\]\[9\] _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__and3_1
X_8710_ reg_data\[19\]\[27\] _3185_ _4274_ vssd1 vssd1 vccd1 vccd1 _4282_ sky130_fd_sc_hd__mux2_1
X_6971_ _3262_ reg_data\[10\]\[29\] _3331_ vssd1 vssd1 vccd1 vccd1 _3341_ sky130_fd_sc_hd__mux2_1
X_5922_ reg_data\[14\]\[23\] _2301_ _1958_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__and3_1
X_9690_ clknet_leaf_1_i_clk _0834_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8641_ _4245_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__clkbuf_1
X_5853_ reg_data\[14\]\[22\] _2301_ _1958_ vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__and3_1
X_8572_ reg_data\[1\]\[26\] _3183_ _4202_ vssd1 vssd1 vccd1 vccd1 _4209_ sky130_fd_sc_hd__mux2_1
X_4804_ reg_data\[16\]\[5\] _1219_ _1221_ reg_data\[9\]\[5\] vssd1 vssd1 vccd1 vccd1
+ _1420_ sky130_fd_sc_hd__a22o_1
X_5784_ reg_data\[24\]\[21\] _1847_ _1848_ reg_data\[28\]\[21\] _2367_ vssd1 vssd1
+ vccd1 vccd1 _2368_ sky130_fd_sc_hd__a221o_1
X_7523_ _3264_ reg_data\[21\]\[30\] _3602_ vssd1 vssd1 vccd1 vccd1 _3636_ sky130_fd_sc_hd__mux2_1
X_4735_ reg_data\[14\]\[4\] _1189_ _1193_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__and3_1
X_7454_ _3598_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__clkbuf_1
X_4666_ reg_data\[5\]\[3\] _1179_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__and3_1
X_7385_ reg_data\[3\]\[30\] _3191_ _3528_ vssd1 vssd1 vccd1 vccd1 _3562_ sky130_fd_sc_hd__mux2_1
X_6405_ reg_data\[17\]\[0\] _2489_ _1395_ vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__and3_1
X_4597_ _1218_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__clkbuf_4
X_6336_ reg_data\[12\]\[31\] _1076_ _1128_ vssd1 vssd1 vccd1 vccd1 _2901_ sky130_fd_sc_hd__and3_1
X_9124_ clknet_leaf_63_i_clk _0268_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_9055_ clknet_leaf_4_i_clk _0199_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6267_ _2834_ vssd1 vssd1 vccd1 vccd1 rdata2\[29\] sky130_fd_sc_hd__clkbuf_1
X_6198_ reg_data\[0\]\[28\] _2427_ _2765_ _2766_ _2767_ vssd1 vssd1 vccd1 vccd1 _2768_
+ sky130_fd_sc_hd__a2111o_1
X_5218_ reg_data\[3\]\[12\] _1815_ _1817_ _1818_ _1819_ vssd1 vssd1 vccd1 vccd1 _1820_
+ sky130_fd_sc_hd__a2111o_1
X_8006_ _3903_ reg_data\[9\]\[21\] _3901_ vssd1 vssd1 vccd1 vccd1 _3904_ sky130_fd_sc_hd__mux2_1
X_5149_ reg_data\[7\]\[11\] _1185_ _1750_ _1751_ _1752_ vssd1 vssd1 vccd1 vccd1 _1753_
+ sky130_fd_sc_hd__a2111o_1
X_8908_ clknet_leaf_28_i_clk _0052_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_9888_ clknet_leaf_38_i_clk _0958_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_8839_ _4350_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__clkbuf_1
X_4520_ _0997_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__clkbuf_4
X_4451_ _1071_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__clkbuf_4
X_7170_ reg_data\[7\]\[25\] _3181_ _3442_ vssd1 vssd1 vccd1 vccd1 _3448_ sky130_fd_sc_hd__mux2_1
X_6121_ reg_data\[7\]\[27\] _2386_ _2691_ _2692_ _2693_ vssd1 vssd1 vccd1 vccd1 _2694_
+ sky130_fd_sc_hd__a2111o_1
X_4382_ i_rs2[0] i_rs2[2] i_rs2[1] i_rs2[3] vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__o31ai_1
X_6052_ reg_data\[22\]\[26\] _2143_ _2256_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__and3_1
X_5003_ reg_data\[23\]\[9\] _1099_ _1101_ reg_data\[19\]\[9\] vssd1 vssd1 vccd1 vccd1
+ _1612_ sky130_fd_sc_hd__a22o_1
X_9811_ clknet_leaf_35_i_clk rdata1\[27\] vssd1 vssd1 vccd1 vccd1 r_data1\[27\] sky130_fd_sc_hd__dfxtp_1
X_9742_ clknet_leaf_23_i_clk _0886_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6954_ _3332_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__clkbuf_1
X_5905_ reg_data\[24\]\[23\] _2409_ _2410_ reg_data\[28\]\[23\] _2485_ vssd1 vssd1
+ vccd1 vccd1 _2486_ sky130_fd_sc_hd__a221o_1
X_9673_ clknet_leaf_44_i_clk _0817_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_8624_ _4236_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__clkbuf_1
X_6885_ reg_data\[2\]\[21\] _3173_ _3293_ vssd1 vssd1 vccd1 vccd1 _3295_ sky130_fd_sc_hd__mux2_1
X_5836_ reg_data\[21\]\[22\] _1883_ _1943_ vssd1 vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__and3_1
X_5767_ reg_data\[3\]\[21\] _1815_ _2348_ _2349_ _2350_ vssd1 vssd1 vccd1 vccd1 _2351_
+ sky130_fd_sc_hd__a2111o_1
X_8555_ reg_data\[1\]\[18\] _3166_ _4191_ vssd1 vssd1 vccd1 vccd1 _4200_ sky130_fd_sc_hd__mux2_1
X_7506_ _3627_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__clkbuf_1
X_8486_ _4163_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__clkbuf_1
X_5698_ _2284_ vssd1 vssd1 vccd1 vccd1 rdata1\[20\] sky130_fd_sc_hd__clkbuf_1
X_4718_ reg_data\[22\]\[4\] _1143_ _1270_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__and3_1
X_7437_ _3248_ reg_data\[20\]\[22\] _3587_ vssd1 vssd1 vccd1 vccd1 _3590_ sky130_fd_sc_hd__mux2_1
X_4649_ _1269_ vssd1 vssd1 vccd1 vccd1 rdata1\[3\] sky130_fd_sc_hd__clkbuf_1
X_7368_ _3553_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__clkbuf_1
X_9107_ clknet_leaf_18_i_clk _0251_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6319_ reg_data\[24\]\[30\] _2453_ _2454_ reg_data\[28\]\[30\] _2884_ vssd1 vssd1
+ vccd1 vccd1 _2885_ sky130_fd_sc_hd__a221o_1
X_7299_ reg_data\[5\]\[21\] _3173_ _3515_ vssd1 vssd1 vccd1 vccd1 _3517_ sky130_fd_sc_hd__mux2_1
X_9038_ clknet_leaf_38_i_clk _0182_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6670_ _3153_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__clkbuf_1
X_5621_ reg_data\[5\]\[19\] _2097_ _1925_ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__and3_1
X_5552_ _1038_ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__clkbuf_4
X_8340_ _4086_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__clkbuf_1
X_4503_ _1062_ _1094_ _1114_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__and3_4
X_8271_ _4049_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__clkbuf_1
X_5483_ reg_data\[1\]\[16\] _1904_ _1905_ reg_data\[15\]\[16\] vssd1 vssd1 vccd1 vccd1
+ _2077_ sky130_fd_sc_hd__a22o_1
X_4434_ reg_data\[30\]\[2\] _1055_ _1056_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__and3_1
X_7222_ _3475_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__clkbuf_1
X_4365_ rs2\[4\] i_rs2[4] _0994_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__mux2_1
X_7153_ reg_data\[7\]\[17\] _3164_ _3431_ vssd1 vssd1 vccd1 vccd1 _3439_ sky130_fd_sc_hd__mux2_1
X_6104_ _2669_ _2673_ _2675_ _2677_ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__or4_1
X_7084_ _3237_ reg_data\[8\]\[17\] _3394_ vssd1 vssd1 vccd1 vccd1 _3402_ sky130_fd_sc_hd__mux2_1
X_6035_ reg_data\[5\]\[25\] _2430_ _1338_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_42_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_7986_ i_data[15] vssd1 vssd1 vccd1 vccd1 _3890_ sky130_fd_sc_hd__clkbuf_4
X_9725_ clknet_leaf_4_i_clk _0869_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6937_ _3323_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__clkbuf_1
X_9656_ clknet_leaf_10_i_clk _0800_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6868_ reg_data\[2\]\[13\] _3156_ _3282_ vssd1 vssd1 vccd1 vccd1 _3286_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_57_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_9587_ clknet_leaf_34_i_clk _0731_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5819_ reg_data\[27\]\[22\] _2392_ _2395_ _2398_ _2401_ vssd1 vssd1 vccd1 vccd1 _2402_
+ sky130_fd_sc_hd__a2111o_1
X_8607_ _3879_ reg_data\[12\]\[10\] _4227_ vssd1 vssd1 vccd1 vccd1 _4228_ sky130_fd_sc_hd__mux2_1
X_6799_ _3242_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__clkbuf_1
X_8538_ _4179_ vssd1 vssd1 vccd1 vccd1 _4191_ sky130_fd_sc_hd__buf_4
X_8469_ _4154_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__clkbuf_1
X_7840_ _3239_ reg_data\[27\]\[18\] _3796_ vssd1 vssd1 vccd1 vccd1 _3805_ sky130_fd_sc_hd__mux2_1
X_7771_ _3768_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__clkbuf_1
X_4983_ reg_data\[17\]\[9\] _1042_ _1238_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__and3_1
X_6722_ _3188_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__clkbuf_1
X_9510_ clknet_leaf_45_i_clk _0654_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_9441_ clknet_leaf_73_i_clk _0585_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6653_ reg_data\[4\]\[6\] _3141_ _3129_ vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__mux2_1
X_5604_ reg_data\[8\]\[18\] _1841_ _1842_ reg_data\[10\]\[18\] _2193_ vssd1 vssd1
+ vccd1 vccd1 _2194_ sky130_fd_sc_hd__a221o_1
X_9372_ clknet_leaf_74_i_clk _0516_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6584_ r_data2\[13\] _3094_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__and2_1
X_5535_ reg_data\[5\]\[17\] _1824_ _1954_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__and3_1
X_8323_ _4077_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__clkbuf_1
X_8254_ _4040_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__clkbuf_1
X_5466_ reg_data\[18\]\[16\] _1816_ _1513_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__and3_1
X_4417_ rs1_mux\[0\] _1026_ _1030_ _1033_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__and4_2
X_7205_ _3466_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__clkbuf_1
X_5397_ reg_data\[27\]\[15\] _1786_ _1991_ _1992_ _1993_ vssd1 vssd1 vccd1 vccd1 _1994_
+ sky130_fd_sc_hd__a2111o_1
X_8185_ _3867_ reg_data\[14\]\[4\] _3999_ vssd1 vssd1 vccd1 vccd1 _4004_ sky130_fd_sc_hd__mux2_1
X_7136_ reg_data\[7\]\[9\] _3147_ _3420_ vssd1 vssd1 vccd1 vccd1 _3430_ sky130_fd_sc_hd__mux2_1
X_7067_ _3220_ reg_data\[8\]\[9\] _3383_ vssd1 vssd1 vccd1 vccd1 _3393_ sky130_fd_sc_hd__mux2_1
X_6018_ reg_data\[27\]\[25\] _2392_ _2592_ _2593_ _2594_ vssd1 vssd1 vccd1 vccd1 _2595_
+ sky130_fd_sc_hd__a2111o_1
X_7969_ _3878_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__clkbuf_1
X_9708_ clknet_leaf_40_i_clk _0852_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_9639_ clknet_leaf_48_i_clk _0783_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_5320_ _1056_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__clkbuf_4
X_5251_ _1832_ _1840_ _1846_ _1852_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__or4_1
X_5182_ _1769_ _1774_ _1779_ _1784_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__or4_1
X_8941_ clknet_leaf_40_i_clk _0085_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_8872_ clknet_leaf_49_i_clk _0016_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_7823_ _3784_ vssd1 vssd1 vccd1 vccd1 _3796_ sky130_fd_sc_hd__buf_4
X_7754_ _3759_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__clkbuf_1
X_6705_ i_data[23] vssd1 vssd1 vccd1 vccd1 _3177_ sky130_fd_sc_hd__clkbuf_4
X_4966_ _1190_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__buf_2
X_7685_ _3220_ reg_data\[25\]\[9\] _3713_ vssd1 vssd1 vccd1 vccd1 _3723_ sky130_fd_sc_hd__mux2_1
X_4897_ _1138_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__buf_2
X_9424_ clknet_leaf_34_i_clk _0568_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6636_ _3130_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__clkbuf_1
X_9355_ clknet_leaf_59_i_clk _0499_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6567_ r_data2\[5\] _3083_ vssd1 vssd1 vccd1 vccd1 _3089_ sky130_fd_sc_hd__and2_1
X_8306_ _4067_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__clkbuf_1
X_5518_ reg_data\[8\]\[17\] _1797_ _1798_ reg_data\[10\]\[17\] _2110_ vssd1 vssd1
+ vccd1 vccd1 _2111_ sky130_fd_sc_hd__a221o_1
X_6498_ r_data1\[5\] _3046_ vssd1 vssd1 vccd1 vccd1 _3052_ sky130_fd_sc_hd__and2_1
X_9286_ clknet_leaf_54_i_clk _0430_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8237_ _3919_ reg_data\[14\]\[29\] _4021_ vssd1 vssd1 vccd1 vccd1 _4031_ sky130_fd_sc_hd__mux2_1
X_5449_ reg_data\[13\]\[16\] _1608_ _1257_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__and3_1
X_8168_ _3994_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__clkbuf_1
X_7119_ _3421_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_1
X_8099_ _3957_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__clkbuf_1
X_4820_ reg_data\[5\]\[6\] _1076_ _1250_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__and3_1
X_4751_ reg_data\[17\]\[5\] _1042_ _1238_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__and3_1
X_4682_ reg_data\[16\]\[3\] _1219_ _1221_ reg_data\[9\]\[3\] vssd1 vssd1 vccd1 vccd1
+ _1302_ sky130_fd_sc_hd__a22o_1
X_7470_ _3608_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__clkbuf_1
X_6421_ reg_data\[23\]\[0\] _1205_ _1208_ reg_data\[19\]\[0\] vssd1 vssd1 vccd1 vccd1
+ _2983_ sky130_fd_sc_hd__a22o_1
X_9140_ clknet_leaf_18_i_clk _0284_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6352_ reg_data\[22\]\[31\] _1207_ _1151_ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__and3_1
X_9071_ clknet_leaf_23_i_clk _0215_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6283_ reg_data\[7\]\[30\] _2386_ _2847_ _2848_ _2849_ vssd1 vssd1 vccd1 vccd1 _2850_
+ sky130_fd_sc_hd__a2111o_1
X_5303_ reg_data\[2\]\[13\] _1837_ _1901_ _1902_ reg_data\[11\]\[13\] vssd1 vssd1
+ vccd1 vccd1 _1903_ sky130_fd_sc_hd__a32o_1
X_8022_ _3914_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__clkbuf_1
X_5234_ reg_data\[23\]\[12\] _1834_ _1835_ reg_data\[19\]\[12\] vssd1 vssd1 vccd1
+ vccd1 _1836_ sky130_fd_sc_hd__a22o_1
X_5165_ reg_data\[21\]\[12\] _1480_ _1240_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__and3_1
X_5096_ reg_data\[16\]\[10\] _1219_ _1221_ reg_data\[9\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _1702_ sky130_fd_sc_hd__a22o_1
X_8924_ clknet_leaf_75_i_clk _0068_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_8855_ _4358_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__clkbuf_1
X_7806_ _3787_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__clkbuf_1
X_5998_ reg_data\[22\]\[25\] _2143_ _2256_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__and3_1
X_8786_ _3923_ reg_data\[29\]\[31\] _4287_ vssd1 vssd1 vccd1 vccd1 _4322_ sky130_fd_sc_hd__mux2_1
X_4949_ reg_data\[26\]\[8\] _1132_ _1134_ reg_data\[29\]\[8\] vssd1 vssd1 vccd1 vccd1
+ _1560_ sky130_fd_sc_hd__a22o_1
X_7737_ _3204_ reg_data\[26\]\[1\] _3749_ vssd1 vssd1 vccd1 vccd1 _3751_ sky130_fd_sc_hd__mux2_1
X_7668_ _3714_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__clkbuf_1
X_6619_ r_data2\[30\] _3082_ vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__and2_1
X_9407_ clknet_leaf_68_i_clk _0551_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_7599_ _3195_ reg_data\[24\]\[0\] _3677_ vssd1 vssd1 vccd1 vccd1 _3678_ sky130_fd_sc_hd__mux2_1
X_9338_ clknet_leaf_60_i_clk _0482_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_9269_ clknet_leaf_36_i_clk _0413_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6970_ _3340_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__clkbuf_1
X_5921_ reg_data\[13\]\[23\] _2183_ _2299_ vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__and3_1
X_8640_ _3913_ reg_data\[12\]\[26\] _4238_ vssd1 vssd1 vccd1 vccd1 _4245_ sky130_fd_sc_hd__mux2_1
X_5852_ reg_data\[13\]\[22\] _2183_ _2299_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__and3_1
X_8571_ _4208_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__clkbuf_1
X_4803_ reg_data\[27\]\[5\] _1199_ _1416_ _1417_ _1418_ vssd1 vssd1 vccd1 vccd1 _1419_
+ sky130_fd_sc_hd__a2111o_1
X_5783_ reg_data\[26\]\[21\] _1849_ _1850_ reg_data\[29\]\[21\] vssd1 vssd1 vccd1
+ vccd1 _2367_ sky130_fd_sc_hd__a22o_1
X_7522_ _3635_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__clkbuf_1
X_4734_ reg_data\[13\]\[4\] _1186_ _1191_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__and3_1
X_7453_ _3264_ reg_data\[20\]\[30\] _3564_ vssd1 vssd1 vccd1 vccd1 _3598_ sky130_fd_sc_hd__mux2_1
X_4665_ _1144_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__clkbuf_4
X_7384_ _3561_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__clkbuf_1
X_4596_ _1207_ _1172_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__and2_4
X_6404_ reg_data\[22\]\[0\] _1207_ _1151_ vssd1 vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__and3_1
X_6335_ reg_data\[14\]\[31\] _1082_ _1090_ vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__and3_1
X_9123_ clknet_leaf_66_i_clk _0267_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_9054_ clknet_leaf_4_i_clk _0198_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6266_ _2825_ _2829_ _2831_ _2833_ vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__or4_1
X_8005_ i_data[21] vssd1 vssd1 vccd1 vccd1 _3903_ sky130_fd_sc_hd__buf_4
X_6197_ reg_data\[5\]\[28\] _2430_ _1338_ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__and3_1
X_5217_ reg_data\[20\]\[12\] _1629_ _1743_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__and3_1
X_5148_ reg_data\[13\]\[11\] _1354_ _1191_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__and3_1
X_5079_ reg_data\[30\]\[10\] _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__and3_1
X_8907_ clknet_leaf_44_i_clk _0051_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_9887_ clknet_leaf_34_i_clk _0957_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_8838_ reg_data\[11\]\[23\] i_data[23] _4346_ vssd1 vssd1 vccd1 vccd1 _4350_ sky130_fd_sc_hd__mux2_1
X_8769_ _4313_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__clkbuf_1
X_4450_ reg_data\[4\]\[2\] _1072_ _1059_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__and3_1
X_4381_ _1010_ vssd1 vssd1 vccd1 vccd1 rs2_mux\[2\] sky130_fd_sc_hd__clkinv_2
X_6120_ reg_data\[13\]\[27\] _2214_ _2102_ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__and3_1
X_6051_ _2626_ vssd1 vssd1 vccd1 vccd1 rdata2\[25\] sky130_fd_sc_hd__clkbuf_1
X_5002_ _1594_ _1599_ _1604_ _1610_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__or4_1
X_9810_ clknet_leaf_33_i_clk rdata1\[26\] vssd1 vssd1 vccd1 vccd1 r_data1\[26\] sky130_fd_sc_hd__dfxtp_1
X_9741_ clknet_leaf_16_i_clk _0885_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6953_ _3243_ reg_data\[10\]\[20\] _3331_ vssd1 vssd1 vccd1 vccd1 _3332_ sky130_fd_sc_hd__mux2_1
X_5904_ reg_data\[26\]\[23\] _2411_ _2412_ reg_data\[29\]\[23\] vssd1 vssd1 vccd1
+ vccd1 _2485_ sky130_fd_sc_hd__a22o_1
X_6884_ _3294_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__clkbuf_1
X_9672_ clknet_leaf_46_i_clk _0816_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_5835_ reg_data\[22\]\[22\] _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__and3_1
X_8623_ _3896_ reg_data\[12\]\[18\] _4227_ vssd1 vssd1 vccd1 vccd1 _4236_ sky130_fd_sc_hd__mux2_1
X_5766_ reg_data\[30\]\[21\] _2234_ _1164_ vssd1 vssd1 vccd1 vccd1 _2350_ sky130_fd_sc_hd__and3_1
X_8554_ _4199_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__clkbuf_1
X_7505_ _3246_ reg_data\[21\]\[21\] _3625_ vssd1 vssd1 vccd1 vccd1 _3627_ sky130_fd_sc_hd__mux2_1
X_8485_ _3894_ reg_data\[18\]\[17\] _4155_ vssd1 vssd1 vccd1 vccd1 _4163_ sky130_fd_sc_hd__mux2_1
X_4717_ _1335_ vssd1 vssd1 vccd1 vccd1 rdata1\[4\] sky130_fd_sc_hd__clkbuf_1
X_5697_ _2275_ _2279_ _2281_ _2283_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__or4_1
X_7436_ _3589_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__clkbuf_1
X_4648_ _1260_ _1264_ _1266_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__or4_1
X_9106_ clknet_leaf_18_i_clk _0250_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_7367_ reg_data\[3\]\[21\] _3173_ _3551_ vssd1 vssd1 vccd1 vccd1 _3553_ sky130_fd_sc_hd__mux2_1
X_4579_ reg_data\[2\]\[2\] _1001_ _1168_ _1200_ reg_data\[11\]\[2\] vssd1 vssd1 vccd1
+ vccd1 _1201_ sky130_fd_sc_hd__a32o_1
X_6318_ reg_data\[26\]\[30\] _2455_ _2456_ reg_data\[29\]\[30\] vssd1 vssd1 vccd1
+ vccd1 _2884_ sky130_fd_sc_hd__a22o_1
X_7298_ _3516_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__clkbuf_1
X_6249_ reg_data\[6\]\[29\] _2555_ _1270_ vssd1 vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__and3_1
X_9037_ clknet_leaf_50_i_clk _0181_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5620_ reg_data\[4\]\[19\] _1718_ _1863_ vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__and3_1
X_5551_ _2142_ vssd1 vssd1 vccd1 vccd1 rdata2\[17\] sky130_fd_sc_hd__clkbuf_1
X_8270_ _3884_ reg_data\[15\]\[12\] _4046_ vssd1 vssd1 vccd1 vccd1 _4049_ sky130_fd_sc_hd__mux2_1
X_4502_ reg_data\[8\]\[2\] _1116_ _1119_ reg_data\[10\]\[2\] _1124_ vssd1 vssd1 vccd1
+ vccd1 _1125_ sky130_fd_sc_hd__a221o_1
X_5482_ reg_data\[2\]\[16\] _1837_ _1901_ _1902_ reg_data\[11\]\[16\] vssd1 vssd1
+ vccd1 vccd1 _2076_ sky130_fd_sc_hd__a32o_1
X_7221_ reg_data\[6\]\[17\] _3164_ _3467_ vssd1 vssd1 vccd1 vccd1 _3475_ sky130_fd_sc_hd__mux2_1
X_4433_ rs1_mux\[0\] _1025_ rs1_mux\[2\] rs1_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1056_
+ sky130_fd_sc_hd__and4bb_2
X_4364_ i_rs2[0] i_rs2[3] i_rs2[2] i_rs2[1] vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__or4_1
X_7152_ _3438_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__clkbuf_1
X_6103_ reg_data\[24\]\[26\] _2453_ _2454_ reg_data\[28\]\[26\] _2676_ vssd1 vssd1
+ vccd1 vccd1 _2677_ sky130_fd_sc_hd__a221o_1
X_7083_ _3401_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_1
X_6034_ reg_data\[4\]\[25\] _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__and3_1
X_7985_ _3889_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__clkbuf_1
X_6936_ _3227_ reg_data\[10\]\[12\] _3320_ vssd1 vssd1 vccd1 vccd1 _3323_ sky130_fd_sc_hd__mux2_1
X_9724_ clknet_leaf_11_i_clk _0868_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_9655_ clknet_leaf_24_i_clk _0799_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6867_ _3285_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__clkbuf_1
X_9586_ clknet_leaf_34_i_clk _0730_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_5818_ reg_data\[1\]\[22\] _2336_ _2399_ _2400_ reg_data\[15\]\[22\] vssd1 vssd1
+ vccd1 vccd1 _2401_ sky130_fd_sc_hd__a32o_1
X_8606_ _4215_ vssd1 vssd1 vccd1 vccd1 _4227_ sky130_fd_sc_hd__buf_4
X_6798_ _3241_ reg_data\[22\]\[19\] _3223_ vssd1 vssd1 vccd1 vccd1 _3242_ sky130_fd_sc_hd__mux2_1
X_8537_ _4190_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__clkbuf_1
X_5749_ reg_data\[23\]\[21\] _1787_ _1788_ reg_data\[19\]\[21\] vssd1 vssd1 vccd1
+ vccd1 _2334_ sky130_fd_sc_hd__a22o_1
X_8468_ _3877_ reg_data\[18\]\[9\] _4144_ vssd1 vssd1 vccd1 vccd1 _4154_ sky130_fd_sc_hd__mux2_1
X_7419_ _3580_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__clkbuf_1
X_8399_ _4117_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__clkbuf_1
X_7770_ _3237_ reg_data\[26\]\[17\] _3760_ vssd1 vssd1 vccd1 vccd1 _3768_ sky130_fd_sc_hd__mux2_1
X_4982_ reg_data\[22\]\[9\] _1536_ _1236_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__and3_1
X_6721_ reg_data\[4\]\[28\] _3187_ _3171_ vssd1 vssd1 vccd1 vccd1 _3188_ sky130_fd_sc_hd__mux2_1
X_6652_ i_data[6] vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__buf_2
X_9440_ clknet_leaf_74_i_clk _0584_ vssd1 vssd1 vccd1 vccd1 reg_data\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_9371_ clknet_leaf_74_i_clk _0515_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5603_ reg_data\[16\]\[18\] _1843_ _1844_ reg_data\[9\]\[18\] vssd1 vssd1 vccd1 vccd1
+ _2193_ sky130_fd_sc_hd__a22o_1
X_8322_ _3867_ reg_data\[16\]\[4\] _4072_ vssd1 vssd1 vccd1 vccd1 _4077_ sky130_fd_sc_hd__mux2_1
X_6583_ _3097_ vssd1 vssd1 vccd1 vccd1 o_data2[12] sky130_fd_sc_hd__buf_2
X_5534_ reg_data\[4\]\[17\] _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__and3_1
X_8253_ _3867_ reg_data\[15\]\[4\] _4035_ vssd1 vssd1 vccd1 vccd1 _4040_ sky130_fd_sc_hd__mux2_1
X_5465_ reg_data\[25\]\[16\] _1810_ _2056_ _2057_ _2058_ vssd1 vssd1 vccd1 vccd1 _2059_
+ sky130_fd_sc_hd__a2111o_1
X_4416_ _1038_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__buf_2
X_7204_ reg_data\[6\]\[9\] _3147_ _3456_ vssd1 vssd1 vccd1 vccd1 _3466_ sky130_fd_sc_hd__mux2_1
X_8184_ _4003_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__clkbuf_1
X_5396_ reg_data\[1\]\[15\] _1729_ _1793_ _1794_ reg_data\[15\]\[15\] vssd1 vssd1
+ vccd1 vccd1 _1993_ sky130_fd_sc_hd__a32o_1
X_7135_ _3429_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
X_7066_ _3392_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
X_6017_ reg_data\[1\]\[25\] _2336_ _2399_ _2400_ reg_data\[15\]\[25\] vssd1 vssd1
+ vccd1 vccd1 _2594_ sky130_fd_sc_hd__a32o_1
X_7968_ _3877_ reg_data\[9\]\[9\] _3859_ vssd1 vssd1 vccd1 vccd1 _3878_ sky130_fd_sc_hd__mux2_1
X_9707_ clknet_leaf_59_i_clk _0851_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6919_ _3210_ reg_data\[10\]\[4\] _3309_ vssd1 vssd1 vccd1 vccd1 _3314_ sky130_fd_sc_hd__mux2_1
X_7899_ _3229_ reg_data\[28\]\[13\] _3833_ vssd1 vssd1 vccd1 vccd1 _3837_ sky130_fd_sc_hd__mux2_1
X_9638_ clknet_leaf_50_i_clk _0782_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_9569_ clknet_leaf_1_i_clk _0713_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_41_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5250_ reg_data\[24\]\[12\] _1847_ _1848_ reg_data\[28\]\[12\] _1851_ vssd1 vssd1
+ vccd1 vccd1 _1852_ sky130_fd_sc_hd__a221o_1
X_5181_ reg_data\[7\]\[12\] _1780_ _1781_ _1782_ _1783_ vssd1 vssd1 vccd1 vccd1 _1784_
+ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_56_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_8940_ clknet_leaf_40_i_clk _0084_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8871_ clknet_leaf_48_i_clk _0015_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_7822_ _3795_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__clkbuf_1
X_4965_ _1171_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__buf_2
X_7753_ _3220_ reg_data\[26\]\[9\] _3749_ vssd1 vssd1 vccd1 vccd1 _3759_ sky130_fd_sc_hd__mux2_1
X_6704_ _3176_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__clkbuf_1
X_9423_ clknet_leaf_34_i_clk _0567_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_7684_ _3722_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__clkbuf_1
X_4896_ reg_data\[17\]\[7\] _1272_ _1148_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__and3_1
X_6635_ reg_data\[4\]\[0\] _3118_ _3129_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__mux2_1
X_9354_ clknet_leaf_53_i_clk _0498_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6566_ _3088_ vssd1 vssd1 vccd1 vccd1 o_data2[4] sky130_fd_sc_hd__buf_2
X_8305_ _3919_ reg_data\[15\]\[29\] _4057_ vssd1 vssd1 vccd1 vccd1 _4067_ sky130_fd_sc_hd__mux2_1
X_9285_ clknet_leaf_52_i_clk _0429_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5517_ reg_data\[16\]\[17\] _1799_ _1800_ reg_data\[9\]\[17\] vssd1 vssd1 vccd1 vccd1
+ _2110_ sky130_fd_sc_hd__a22o_1
X_8236_ _4030_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__clkbuf_1
X_6497_ _3051_ vssd1 vssd1 vccd1 vccd1 o_data1[4] sky130_fd_sc_hd__buf_2
X_5448_ reg_data\[12\]\[16\] _1986_ _1606_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__and3_1
X_8167_ _3917_ reg_data\[13\]\[28\] _3985_ vssd1 vssd1 vccd1 vccd1 _3994_ sky130_fd_sc_hd__mux2_1
X_5379_ reg_data\[25\]\[15\] _1764_ _1973_ _1974_ _1975_ vssd1 vssd1 vccd1 vccd1 _1976_
+ sky130_fd_sc_hd__a2111o_1
X_8098_ _3917_ reg_data\[30\]\[28\] _3948_ vssd1 vssd1 vccd1 vccd1 _3957_ sky130_fd_sc_hd__mux2_1
X_7118_ reg_data\[7\]\[0\] _3118_ _3420_ vssd1 vssd1 vccd1 vccd1 _3421_ sky130_fd_sc_hd__mux2_1
X_7049_ _3195_ reg_data\[8\]\[0\] _3383_ vssd1 vssd1 vccd1 vccd1 _3384_ sky130_fd_sc_hd__mux2_1
X_4750_ reg_data\[22\]\[5\] _1039_ _1236_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__and3_1
X_4681_ reg_data\[27\]\[3\] _1199_ _1294_ _1297_ _1300_ vssd1 vssd1 vccd1 vccd1 _1301_
+ sky130_fd_sc_hd__a2111o_1
X_6420_ _2969_ _2973_ _2977_ _2981_ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__or4_2
X_6351_ reg_data\[25\]\[31\] _1207_ _1139_ vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__and3_1
X_5302_ _1200_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__clkbuf_4
X_9070_ clknet_leaf_29_i_clk _0214_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6282_ reg_data\[14\]\[30\] _1076_ _1090_ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__and3_1
X_8021_ _3913_ reg_data\[9\]\[26\] _3901_ vssd1 vssd1 vccd1 vccd1 _3914_ sky130_fd_sc_hd__mux2_1
X_5233_ _1208_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__clkbuf_4
X_5164_ reg_data\[17\]\[12\] _1766_ _1708_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__and3_1
X_5095_ reg_data\[27\]\[10\] _1199_ _1698_ _1699_ _1700_ vssd1 vssd1 vccd1 vccd1 _1701_
+ sky130_fd_sc_hd__a2111o_1
X_8923_ clknet_leaf_75_i_clk _0067_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_8854_ reg_data\[11\]\[31\] i_data[31] _4323_ vssd1 vssd1 vccd1 vccd1 _4358_ sky130_fd_sc_hd__mux2_1
X_7805_ _3204_ reg_data\[27\]\[1\] _3785_ vssd1 vssd1 vccd1 vccd1 _3787_ sky130_fd_sc_hd__mux2_1
X_5997_ _2574_ vssd1 vssd1 vccd1 vccd1 rdata2\[24\] sky130_fd_sc_hd__clkbuf_1
X_8785_ _4321_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__clkbuf_1
X_7736_ _3750_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__clkbuf_1
X_4948_ reg_data\[8\]\[8\] _1116_ _1119_ reg_data\[10\]\[8\] _1558_ vssd1 vssd1 vccd1
+ vccd1 _1559_ sky130_fd_sc_hd__a221o_1
X_7667_ _3195_ reg_data\[25\]\[0\] _3713_ vssd1 vssd1 vccd1 vccd1 _3714_ sky130_fd_sc_hd__mux2_1
X_4879_ reg_data\[0\]\[7\] _1070_ _1488_ _1489_ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_
+ sky130_fd_sc_hd__a2111o_1
X_6618_ _3115_ vssd1 vssd1 vccd1 vccd1 o_data2[29] sky130_fd_sc_hd__buf_2
X_9406_ clknet_leaf_71_i_clk _0550_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_7598_ _3676_ vssd1 vssd1 vccd1 vccd1 _3677_ sky130_fd_sc_hd__buf_4
X_9337_ clknet_leaf_67_i_clk _0481_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6549_ _3078_ vssd1 vssd1 vccd1 vccd1 o_data1[29] sky130_fd_sc_hd__buf_2
X_9268_ clknet_leaf_36_i_clk _0412_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_9199_ clknet_leaf_30_i_clk _0343_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_8219_ _3900_ reg_data\[14\]\[20\] _4021_ vssd1 vssd1 vccd1 vccd1 _4022_ sky130_fd_sc_hd__mux2_1
X_5920_ reg_data\[0\]\[23\] _2427_ _2497_ _2498_ _2499_ vssd1 vssd1 vccd1 vccd1 _2500_
+ sky130_fd_sc_hd__a2111o_1
X_5851_ _1184_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__clkbuf_4
X_8570_ reg_data\[1\]\[25\] _3181_ _4202_ vssd1 vssd1 vccd1 vccd1 _4208_ sky130_fd_sc_hd__mux2_1
X_4802_ reg_data\[1\]\[5\] _1298_ _1299_ reg_data\[15\]\[5\] vssd1 vssd1 vccd1 vccd1
+ _1418_ sky130_fd_sc_hd__a22o_1
X_5782_ reg_data\[8\]\[21\] _1841_ _1842_ reg_data\[10\]\[21\] _2365_ vssd1 vssd1
+ vccd1 vccd1 _2366_ sky130_fd_sc_hd__a221o_1
X_7521_ _3262_ reg_data\[21\]\[29\] _3625_ vssd1 vssd1 vccd1 vccd1 _3635_ sky130_fd_sc_hd__mux2_1
X_4733_ reg_data\[0\]\[4\] _1174_ _1348_ _1349_ _1350_ vssd1 vssd1 vccd1 vccd1 _1351_
+ sky130_fd_sc_hd__a2111o_1
X_7452_ _3597_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__clkbuf_1
X_6403_ _2965_ vssd1 vssd1 vccd1 vccd1 rdata1\[0\] sky130_fd_sc_hd__clkbuf_1
X_4664_ reg_data\[4\]\[3\] _1177_ _1283_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__and3_1
X_7383_ reg_data\[3\]\[29\] _3189_ _3551_ vssd1 vssd1 vccd1 vccd1 _3561_ sky130_fd_sc_hd__mux2_1
X_4595_ _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__clkbuf_4
X_6334_ reg_data\[13\]\[31\] _2473_ _1086_ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__and3_1
X_9122_ clknet_leaf_66_i_clk _0266_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6265_ reg_data\[24\]\[29\] _2453_ _2454_ reg_data\[28\]\[29\] _2832_ vssd1 vssd1
+ vccd1 vccd1 _2833_ sky130_fd_sc_hd__a221o_1
X_9053_ clknet_leaf_4_i_clk _0197_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_5216_ reg_data\[30\]\[12\] _1401_ _1402_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__and3_1
X_8004_ _3902_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__clkbuf_1
X_6196_ reg_data\[4\]\[28\] _1175_ _1342_ vssd1 vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__and3_1
X_5147_ reg_data\[12\]\[11\] _1693_ _1289_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__and3_1
X_5078_ reg_data\[18\]\[10\] _1159_ _1513_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__and3_1
X_8906_ clknet_leaf_40_i_clk _0050_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_9886_ clknet_leaf_31_i_clk _0956_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_8837_ _4349_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__clkbuf_1
X_8768_ _3905_ reg_data\[29\]\[22\] _4310_ vssd1 vssd1 vccd1 vccd1 _4313_ sky130_fd_sc_hd__mux2_1
X_7719_ _3254_ reg_data\[25\]\[25\] _3735_ vssd1 vssd1 vccd1 vccd1 _3741_ sky130_fd_sc_hd__mux2_1
X_8699_ _4276_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__clkbuf_1
X_4380_ _0994_ _1007_ _1008_ _1009_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__a31o_2
X_6050_ _2617_ _2621_ _2623_ _2625_ vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__or4_1
X_5001_ reg_data\[7\]\[9\] _1081_ _1605_ _1607_ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_
+ sky130_fd_sc_hd__a2111o_1
X_9740_ clknet_leaf_23_i_clk _0884_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6952_ _3308_ vssd1 vssd1 vccd1 vccd1 _3331_ sky130_fd_sc_hd__buf_4
X_5903_ reg_data\[8\]\[23\] _2403_ _2404_ reg_data\[10\]\[23\] _2483_ vssd1 vssd1
+ vccd1 vccd1 _2484_ sky130_fd_sc_hd__a221o_1
X_6883_ reg_data\[2\]\[20\] _3170_ _3293_ vssd1 vssd1 vccd1 vccd1 _3294_ sky130_fd_sc_hd__mux2_1
X_9671_ clknet_leaf_47_i_clk _0815_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_5834_ _1140_ vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__clkbuf_4
X_8622_ _4235_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__clkbuf_1
X_5765_ reg_data\[20\]\[21\] _2005_ _1160_ vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__and3_1
X_8553_ reg_data\[1\]\[17\] _3164_ _4191_ vssd1 vssd1 vccd1 vccd1 _4199_ sky130_fd_sc_hd__mux2_1
X_7504_ _3626_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_3__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4716_ _1326_ _1330_ _1332_ _1334_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__or4_1
X_5696_ reg_data\[24\]\[20\] _1803_ _1804_ reg_data\[28\]\[20\] _2282_ vssd1 vssd1
+ vccd1 vccd1 _2283_ sky130_fd_sc_hd__a221o_1
X_8484_ _4162_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__clkbuf_1
X_7435_ _3246_ reg_data\[20\]\[21\] _3587_ vssd1 vssd1 vccd1 vccd1 _3589_ sky130_fd_sc_hd__mux2_1
X_4647_ reg_data\[24\]\[3\] _1127_ _1130_ reg_data\[28\]\[3\] _1267_ vssd1 vssd1 vccd1
+ vccd1 _1268_ sky130_fd_sc_hd__a221o_1
X_7366_ _3552_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__clkbuf_1
X_9105_ clknet_leaf_21_i_clk _0249_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6317_ reg_data\[8\]\[30\] _2447_ _2448_ reg_data\[10\]\[30\] _2882_ vssd1 vssd1
+ vccd1 vccd1 _2883_ sky130_fd_sc_hd__a221o_1
X_4578_ _1000_ _1197_ _1156_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__and3_4
X_7297_ reg_data\[5\]\[20\] _3170_ _3515_ vssd1 vssd1 vccd1 vccd1 _3516_ sky130_fd_sc_hd__mux2_1
X_6248_ reg_data\[3\]\[29\] _2421_ _2813_ _2814_ _2815_ vssd1 vssd1 vccd1 vccd1 _2816_
+ sky130_fd_sc_hd__a2111o_1
X_9036_ clknet_leaf_50_i_clk _0180_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6179_ reg_data\[1\]\[28\] _2336_ _2399_ _2400_ reg_data\[15\]\[28\] vssd1 vssd1
+ vccd1 vccd1 _2750_ sky130_fd_sc_hd__a32o_1
X_9869_ clknet_leaf_61_i_clk _0939_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_5550_ _2133_ _2137_ _2139_ _2141_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__or4_1
X_4501_ reg_data\[16\]\[2\] _1121_ _1123_ reg_data\[9\]\[2\] vssd1 vssd1 vccd1 vccd1
+ _1124_ sky130_fd_sc_hd__a22o_1
X_5481_ reg_data\[23\]\[16\] _1834_ _1835_ reg_data\[19\]\[16\] vssd1 vssd1 vccd1
+ vccd1 _2075_ sky130_fd_sc_hd__a22o_1
X_7220_ _3474_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__clkbuf_1
X_4432_ _1038_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__buf_2
X_4363_ _0994_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__inv_2
X_7151_ reg_data\[7\]\[16\] _3162_ _3431_ vssd1 vssd1 vccd1 vccd1 _3438_ sky130_fd_sc_hd__mux2_1
X_6102_ reg_data\[26\]\[26\] _2455_ _2456_ reg_data\[29\]\[26\] vssd1 vssd1 vccd1
+ vccd1 _2676_ sky130_fd_sc_hd__a22o_1
X_7082_ _3235_ reg_data\[8\]\[16\] _3394_ vssd1 vssd1 vccd1 vccd1 _3401_ sky130_fd_sc_hd__mux2_1
X_6033_ reg_data\[6\]\[25\] _2555_ _2237_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__and3_1
X_7984_ _3888_ reg_data\[9\]\[14\] _3880_ vssd1 vssd1 vccd1 vccd1 _3889_ sky130_fd_sc_hd__mux2_1
X_6935_ _3322_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__clkbuf_1
X_9723_ clknet_leaf_4_i_clk _0867_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_9654_ clknet_leaf_23_i_clk _0798_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6866_ reg_data\[2\]\[12\] _3154_ _3282_ vssd1 vssd1 vccd1 vccd1 _3285_ sky130_fd_sc_hd__mux2_1
X_9585_ clknet_leaf_34_i_clk _0729_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_5817_ _1110_ vssd1 vssd1 vccd1 vccd1 _2400_ sky130_fd_sc_hd__clkbuf_4
X_6797_ i_data[19] vssd1 vssd1 vccd1 vccd1 _3241_ sky130_fd_sc_hd__buf_2
X_8605_ _4226_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__clkbuf_1
X_5748_ _2318_ _2322_ _2328_ _2332_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__or4_2
X_8536_ reg_data\[1\]\[9\] _3147_ _4180_ vssd1 vssd1 vccd1 vccd1 _4190_ sky130_fd_sc_hd__mux2_1
X_5679_ reg_data\[6\]\[20\] _2207_ _1716_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__and3_1
X_8467_ _4153_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__clkbuf_1
X_7418_ _3229_ reg_data\[20\]\[13\] _3576_ vssd1 vssd1 vccd1 vccd1 _3580_ sky130_fd_sc_hd__mux2_1
X_8398_ _3875_ reg_data\[17\]\[8\] _4108_ vssd1 vssd1 vccd1 vccd1 _4117_ sky130_fd_sc_hd__mux2_1
X_7349_ _3543_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__clkbuf_1
X_9019_ clknet_leaf_71_i_clk _0163_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_4981_ _1590_ vssd1 vssd1 vccd1 vccd1 rdata2\[8\] sky130_fd_sc_hd__clkbuf_1
X_6720_ i_data[28] vssd1 vssd1 vccd1 vccd1 _3187_ sky130_fd_sc_hd__buf_4
X_6651_ _3140_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__clkbuf_1
X_9370_ clknet_leaf_74_i_clk _0514_ vssd1 vssd1 vccd1 vccd1 reg_data\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_5602_ reg_data\[27\]\[18\] _1833_ _2189_ _2190_ _2191_ vssd1 vssd1 vccd1 vccd1 _2192_
+ sky130_fd_sc_hd__a2111o_1
X_6582_ r_data2\[12\] _3094_ vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__and2_1
X_5533_ reg_data\[6\]\[17\] _1951_ _1632_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__and3_1
X_8321_ _4076_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__clkbuf_1
X_8252_ _4039_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__clkbuf_1
X_5464_ reg_data\[17\]\[16\] _1509_ _1275_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__and3_1
X_4415_ _1017_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__clkbuf_4
X_5395_ reg_data\[2\]\[15\] _1613_ _1790_ _1791_ reg_data\[11\]\[15\] vssd1 vssd1
+ vccd1 vccd1 _1992_ sky130_fd_sc_hd__a32o_1
X_7203_ _3465_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_1
X_8183_ _3865_ reg_data\[14\]\[3\] _3999_ vssd1 vssd1 vccd1 vccd1 _4003_ sky130_fd_sc_hd__mux2_1
X_7134_ reg_data\[7\]\[8\] _3145_ _3420_ vssd1 vssd1 vccd1 vccd1 _3429_ sky130_fd_sc_hd__mux2_1
X_7065_ _3218_ reg_data\[8\]\[8\] _3383_ vssd1 vssd1 vccd1 vccd1 _3392_ sky130_fd_sc_hd__mux2_1
X_6016_ reg_data\[2\]\[25\] _2219_ _2396_ _2397_ reg_data\[11\]\[25\] vssd1 vssd1
+ vccd1 vccd1 _2593_ sky130_fd_sc_hd__a32o_1
X_7967_ i_data[9] vssd1 vssd1 vccd1 vccd1 _3877_ sky130_fd_sc_hd__buf_2
X_9706_ clknet_leaf_56_i_clk _0850_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6918_ _3313_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__clkbuf_1
X_7898_ _3836_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__clkbuf_1
X_6849_ reg_data\[2\]\[4\] _3137_ _3271_ vssd1 vssd1 vccd1 vccd1 _3276_ sky130_fd_sc_hd__mux2_1
X_9637_ clknet_leaf_45_i_clk _0781_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_9568_ clknet_leaf_76_i_clk _0712_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8519_ _4181_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__clkbuf_1
X_9499_ clknet_leaf_4_i_clk _0643_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5180_ reg_data\[13\]\[12\] _1608_ _1257_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__and3_1
X_8870_ clknet_leaf_48_i_clk _0014_ vssd1 vssd1 vccd1 vccd1 reg_data\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_7821_ _3220_ reg_data\[27\]\[9\] _3785_ vssd1 vssd1 vccd1 vccd1 _3795_ sky130_fd_sc_hd__mux2_1
X_7752_ _3758_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__clkbuf_1
X_4964_ reg_data\[0\]\[8\] _1174_ _1571_ _1572_ _1573_ vssd1 vssd1 vccd1 vccd1 _1574_
+ sky130_fd_sc_hd__a2111o_1
X_6703_ reg_data\[4\]\[22\] _3175_ _3171_ vssd1 vssd1 vccd1 vccd1 _3176_ sky130_fd_sc_hd__mux2_1
X_9422_ clknet_leaf_39_i_clk _0566_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_7683_ _3218_ reg_data\[25\]\[8\] _3713_ vssd1 vssd1 vccd1 vccd1 _3722_ sky130_fd_sc_hd__mux2_1
X_4895_ reg_data\[22\]\[7\] _1143_ _1270_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__and3_1
X_6634_ _3128_ vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__buf_4
X_9353_ clknet_leaf_58_i_clk _0497_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6565_ r_data2\[4\] _3083_ vssd1 vssd1 vccd1 vccd1 _3088_ sky130_fd_sc_hd__and2_1
X_8304_ _4066_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__clkbuf_1
X_5516_ reg_data\[27\]\[17\] _1786_ _2106_ _2107_ _2108_ vssd1 vssd1 vccd1 vccd1 _2109_
+ sky130_fd_sc_hd__a2111o_1
X_6496_ r_data1\[4\] _3046_ vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__and2_1
X_9284_ clknet_leaf_59_i_clk _0428_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8235_ _3917_ reg_data\[14\]\[28\] _4021_ vssd1 vssd1 vccd1 vccd1 _4030_ sky130_fd_sc_hd__mux2_1
X_5447_ reg_data\[14\]\[16\] _1867_ _1379_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__and3_1
X_8166_ _3993_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__clkbuf_1
X_5378_ reg_data\[21\]\[15\] _1480_ _1240_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__and3_1
X_8097_ _3956_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__clkbuf_1
X_7117_ _3419_ vssd1 vssd1 vccd1 vccd1 _3420_ sky130_fd_sc_hd__buf_4
X_7048_ _3382_ vssd1 vssd1 vccd1 vccd1 _3383_ sky130_fd_sc_hd__buf_4
X_8999_ clknet_leaf_48_i_clk _0143_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_4680_ reg_data\[1\]\[3\] _1298_ _1299_ reg_data\[15\]\[3\] vssd1 vssd1 vccd1 vccd1
+ _1300_ sky130_fd_sc_hd__a22o_1
X_6350_ reg_data\[21\]\[31\] _1207_ _1144_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__and3_1
X_5301_ _1168_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__buf_4
X_6281_ reg_data\[12\]\[30\] _1082_ _2271_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__and3_1
X_8020_ i_data[26] vssd1 vssd1 vccd1 vccd1 _3913_ sky130_fd_sc_hd__clkbuf_4
X_5232_ _1205_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__buf_4
X_5163_ _1038_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__clkbuf_4
X_5094_ reg_data\[1\]\[10\] _1298_ _1299_ reg_data\[15\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _1700_ sky130_fd_sc_hd__a22o_1
X_8922_ clknet_leaf_75_i_clk _0066_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8853_ _4357_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__clkbuf_1
X_7804_ _3786_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__clkbuf_1
X_5996_ _2565_ _2569_ _2571_ _2573_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__or4_1
X_8784_ _3921_ reg_data\[29\]\[30\] _4287_ vssd1 vssd1 vccd1 vccd1 _4321_ sky130_fd_sc_hd__mux2_1
X_7735_ _3195_ reg_data\[26\]\[0\] _3749_ vssd1 vssd1 vccd1 vccd1 _3750_ sky130_fd_sc_hd__mux2_1
X_4947_ reg_data\[16\]\[8\] _1121_ _1123_ reg_data\[9\]\[8\] vssd1 vssd1 vccd1 vccd1
+ _1558_ sky130_fd_sc_hd__a22o_1
X_7666_ _3712_ vssd1 vssd1 vccd1 vccd1 _3713_ sky130_fd_sc_hd__buf_4
X_4878_ reg_data\[4\]\[7\] _1490_ _1315_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__and3_1
X_6617_ r_data2\[29\] _3105_ vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__and2_1
X_9405_ clknet_leaf_69_i_clk _0549_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_7597_ _3381_ _3675_ vssd1 vssd1 vccd1 vccd1 _3676_ sky130_fd_sc_hd__nand2_4
X_9336_ clknet_leaf_69_i_clk _0480_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6548_ r_data1\[29\] _3068_ vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__and2_1
X_9267_ clknet_leaf_36_i_clk _0411_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6479_ reg_data\[16\]\[1\] _1218_ _1220_ reg_data\[9\]\[1\] vssd1 vssd1 vccd1 vccd1
+ _3039_ sky130_fd_sc_hd__a22o_1
X_9198_ clknet_leaf_31_i_clk _0342_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_8218_ _3998_ vssd1 vssd1 vccd1 vccd1 _4021_ sky130_fd_sc_hd__buf_4
X_8149_ _3984_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_40_i_clk clknet_3_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_55_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5850_ reg_data\[0\]\[22\] _2427_ _2428_ _2429_ _2431_ vssd1 vssd1 vccd1 vccd1 _2432_
+ sky130_fd_sc_hd__a2111o_1
X_4801_ reg_data\[2\]\[5\] _1002_ _1295_ _1296_ reg_data\[11\]\[5\] vssd1 vssd1 vccd1
+ vccd1 _1417_ sky130_fd_sc_hd__a32o_1
X_5781_ reg_data\[16\]\[21\] _1843_ _1844_ reg_data\[9\]\[21\] vssd1 vssd1 vccd1 vccd1
+ _2365_ sky130_fd_sc_hd__a22o_1
X_7520_ _3634_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__clkbuf_1
X_4732_ reg_data\[5\]\[4\] _1179_ _1285_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__and3_1
X_4663_ _1160_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__clkbuf_4
X_7451_ _3262_ reg_data\[20\]\[29\] _3587_ vssd1 vssd1 vccd1 vccd1 _3597_ sky130_fd_sc_hd__mux2_1
X_6402_ _2956_ _2960_ _2962_ _2964_ vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__or4_2
X_7382_ _3560_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__clkbuf_1
X_4594_ _1001_ _1215_ _1197_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__and3_4
X_6333_ reg_data\[0\]\[31\] _2381_ _2895_ _2896_ _2897_ vssd1 vssd1 vccd1 vccd1 _2898_
+ sky130_fd_sc_hd__a2111o_1
X_9121_ clknet_leaf_2_i_clk _0265_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6264_ reg_data\[26\]\[29\] _2455_ _2456_ reg_data\[29\]\[29\] vssd1 vssd1 vccd1
+ vccd1 _2832_ sky130_fd_sc_hd__a22o_1
X_9052_ clknet_leaf_12_i_clk _0196_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_5215_ reg_data\[18\]\[12\] _1816_ _1513_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__and3_1
X_8003_ _3900_ reg_data\[9\]\[20\] _3901_ vssd1 vssd1 vccd1 vccd1 _3902_ sky130_fd_sc_hd__mux2_1
X_6195_ reg_data\[6\]\[28\] _2555_ _2237_ vssd1 vssd1 vccd1 vccd1 _2765_ sky130_fd_sc_hd__and3_1
X_5146_ reg_data\[14\]\[11\] _1575_ _1164_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__and3_1
X_5077_ reg_data\[25\]\[10\] _1141_ _1680_ _1681_ _1682_ vssd1 vssd1 vccd1 vccd1 _1683_
+ sky130_fd_sc_hd__a2111o_1
X_8905_ clknet_leaf_49_i_clk _0049_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_9885_ clknet_leaf_35_i_clk _0955_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_8836_ reg_data\[11\]\[22\] i_data[22] _4346_ vssd1 vssd1 vccd1 vccd1 _4349_ sky130_fd_sc_hd__mux2_1
X_5979_ reg_data\[4\]\[24\] _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__and3_1
X_8767_ _4312_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__clkbuf_1
X_7718_ _3740_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__clkbuf_1
X_8698_ reg_data\[19\]\[21\] _3173_ _4274_ vssd1 vssd1 vccd1 vccd1 _4276_ sky130_fd_sc_hd__mux2_1
X_7649_ _3252_ reg_data\[24\]\[24\] _3699_ vssd1 vssd1 vccd1 vccd1 _3704_ sky130_fd_sc_hd__mux2_1
X_9319_ clknet_leaf_48_i_clk _0463_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_5000_ reg_data\[13\]\[9\] _1608_ _1257_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__and3_1
X_6951_ _3330_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__clkbuf_1
X_5902_ reg_data\[16\]\[23\] _2405_ _2406_ reg_data\[9\]\[23\] vssd1 vssd1 vccd1 vccd1
+ _2483_ sky130_fd_sc_hd__a22o_1
X_6882_ _3270_ vssd1 vssd1 vccd1 vccd1 _3293_ sky130_fd_sc_hd__buf_4
X_9670_ clknet_leaf_47_i_clk _0814_ vssd1 vssd1 vccd1 vccd1 reg_data\[18\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_5833_ _2415_ vssd1 vssd1 vccd1 vccd1 rdata1\[22\] sky130_fd_sc_hd__clkbuf_1
X_8621_ _3894_ reg_data\[12\]\[17\] _4227_ vssd1 vssd1 vccd1 vccd1 _4235_ sky130_fd_sc_hd__mux2_1
X_8552_ _4198_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__clkbuf_1
X_7503_ _3243_ reg_data\[21\]\[20\] _3625_ vssd1 vssd1 vccd1 vccd1 _3626_ sky130_fd_sc_hd__mux2_1
X_5764_ reg_data\[18\]\[21\] _1816_ _2120_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__and3_1
X_4715_ reg_data\[24\]\[4\] _1127_ _1130_ reg_data\[28\]\[4\] _1333_ vssd1 vssd1 vccd1
+ vccd1 _1334_ sky130_fd_sc_hd__a221o_1
X_5695_ reg_data\[26\]\[20\] _1805_ _1806_ reg_data\[29\]\[20\] vssd1 vssd1 vccd1
+ vccd1 _2282_ sky130_fd_sc_hd__a22o_1
X_8483_ _3892_ reg_data\[18\]\[16\] _4155_ vssd1 vssd1 vccd1 vccd1 _4162_ sky130_fd_sc_hd__mux2_1
X_7434_ _3588_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__clkbuf_1
X_4646_ reg_data\[26\]\[3\] _1132_ _1134_ reg_data\[29\]\[3\] vssd1 vssd1 vccd1 vccd1
+ _1267_ sky130_fd_sc_hd__a22o_1
X_7365_ reg_data\[3\]\[20\] _3170_ _3551_ vssd1 vssd1 vccd1 vccd1 _3552_ sky130_fd_sc_hd__mux2_1
X_4577_ _1198_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__buf_4
X_9104_ clknet_leaf_23_i_clk _0248_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6316_ reg_data\[16\]\[30\] _2449_ _2450_ reg_data\[9\]\[30\] vssd1 vssd1 vccd1 vccd1
+ _2882_ sky130_fd_sc_hd__a22o_1
X_7296_ _3492_ vssd1 vssd1 vccd1 vccd1 _3515_ sky130_fd_sc_hd__buf_4
X_6247_ reg_data\[30\]\[29\] _1150_ _1164_ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__and3_1
X_9035_ clknet_leaf_52_i_clk _0179_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6178_ reg_data\[2\]\[28\] _2219_ _2396_ _2397_ reg_data\[11\]\[28\] vssd1 vssd1
+ vccd1 vccd1 _2749_ sky130_fd_sc_hd__a32o_1
X_5129_ reg_data\[26\]\[11\] _1132_ _1134_ reg_data\[29\]\[11\] vssd1 vssd1 vccd1
+ vccd1 _1734_ sky130_fd_sc_hd__a22o_1
X_9868_ clknet_leaf_61_i_clk _0938_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8819_ reg_data\[11\]\[14\] i_data[14] _4335_ vssd1 vssd1 vccd1 vccd1 _4340_ sky130_fd_sc_hd__mux2_1
X_9799_ clknet_leaf_54_i_clk rdata1\[15\] vssd1 vssd1 vccd1 vccd1 r_data1\[15\] sky130_fd_sc_hd__dfxtp_1
X_4500_ _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__clkbuf_4
X_5480_ _2059_ _2063_ _2069_ _2073_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__or4_1
X_4431_ _1053_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__clkbuf_4
X_4362_ i_rs_valid vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__buf_2
X_7150_ _3437_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__clkbuf_1
X_6101_ reg_data\[8\]\[26\] _2447_ _2448_ reg_data\[10\]\[26\] _2674_ vssd1 vssd1
+ vccd1 vccd1 _2675_ sky130_fd_sc_hd__a221o_1
X_7081_ _3400_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__clkbuf_1
X_6032_ reg_data\[3\]\[25\] _2421_ _2605_ _2606_ _2607_ vssd1 vssd1 vccd1 vccd1 _2608_
+ sky130_fd_sc_hd__a2111o_1
X_7983_ i_data[14] vssd1 vssd1 vccd1 vccd1 _3888_ sky130_fd_sc_hd__clkbuf_4
X_9722_ clknet_leaf_11_i_clk _0866_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6934_ _3225_ reg_data\[10\]\[11\] _3320_ vssd1 vssd1 vccd1 vccd1 _3322_ sky130_fd_sc_hd__mux2_1
X_9653_ clknet_leaf_20_i_clk _0797_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6865_ _3284_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__clkbuf_1
X_8604_ _3877_ reg_data\[12\]\[9\] _4216_ vssd1 vssd1 vccd1 vccd1 _4226_ sky130_fd_sc_hd__mux2_1
X_9584_ clknet_leaf_34_i_clk _0728_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_5816_ _1108_ vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__clkbuf_4
X_6796_ _3240_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__clkbuf_1
X_5747_ reg_data\[7\]\[21\] _1780_ _2329_ _2330_ _2331_ vssd1 vssd1 vccd1 vccd1 _2332_
+ sky130_fd_sc_hd__a2111o_1
X_8535_ _4189_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__clkbuf_1
X_8466_ _3875_ reg_data\[18\]\[8\] _4144_ vssd1 vssd1 vccd1 vccd1 _4153_ sky130_fd_sc_hd__mux2_1
X_5678_ reg_data\[3\]\[20\] _1770_ _2262_ _2263_ _2264_ vssd1 vssd1 vccd1 vccd1 _2265_
+ sky130_fd_sc_hd__a2111o_1
X_7417_ _3579_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__clkbuf_1
X_8397_ _4116_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__clkbuf_1
X_4629_ _1043_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__clkbuf_4
X_7348_ reg_data\[3\]\[12\] _3154_ _3540_ vssd1 vssd1 vccd1 vccd1 _3543_ sky130_fd_sc_hd__mux2_1
X_7279_ _3506_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__clkbuf_1
X_9018_ clknet_leaf_70_i_clk _0162_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_4980_ _1581_ _1585_ _1587_ _1589_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__or4_4
X_6650_ reg_data\[4\]\[5\] _3139_ _3129_ vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__mux2_1
X_5601_ reg_data\[1\]\[18\] _1904_ _1905_ reg_data\[15\]\[18\] vssd1 vssd1 vccd1 vccd1
+ _2191_ sky130_fd_sc_hd__a22o_1
X_6581_ _3096_ vssd1 vssd1 vccd1 vccd1 o_data2[11] sky130_fd_sc_hd__buf_2
X_8320_ _3865_ reg_data\[16\]\[3\] _4072_ vssd1 vssd1 vccd1 vccd1 _4076_ sky130_fd_sc_hd__mux2_1
X_5532_ reg_data\[3\]\[17\] _1815_ _2121_ _2122_ _2123_ vssd1 vssd1 vccd1 vccd1 _2124_
+ sky130_fd_sc_hd__a2111o_1
X_8251_ _3865_ reg_data\[15\]\[3\] _4035_ vssd1 vssd1 vccd1 vccd1 _4039_ sky130_fd_sc_hd__mux2_1
X_5463_ reg_data\[21\]\[16\] _1883_ _1943_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__and3_1
X_4414_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__clkbuf_4
X_8182_ _4002_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__clkbuf_1
X_5394_ reg_data\[23\]\[15\] _1787_ _1788_ reg_data\[19\]\[15\] vssd1 vssd1 vccd1
+ vccd1 _1991_ sky130_fd_sc_hd__a22o_1
X_7202_ reg_data\[6\]\[8\] _3145_ _3456_ vssd1 vssd1 vccd1 vccd1 _3465_ sky130_fd_sc_hd__mux2_1
X_7133_ _3428_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__clkbuf_1
X_7064_ _3391_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
X_6015_ reg_data\[23\]\[25\] _2393_ _2394_ reg_data\[19\]\[25\] vssd1 vssd1 vccd1
+ vccd1 _2592_ sky130_fd_sc_hd__a22o_1
X_9705_ clknet_leaf_59_i_clk _0849_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_7966_ _3876_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__clkbuf_1
X_6917_ _3208_ reg_data\[10\]\[3\] _3309_ vssd1 vssd1 vccd1 vccd1 _3313_ sky130_fd_sc_hd__mux2_1
X_7897_ _3227_ reg_data\[28\]\[12\] _3833_ vssd1 vssd1 vccd1 vccd1 _3836_ sky130_fd_sc_hd__mux2_1
X_6848_ _3275_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__clkbuf_1
X_9636_ clknet_leaf_47_i_clk _0780_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_9567_ clknet_leaf_0_i_clk _0711_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6779_ i_data[13] vssd1 vssd1 vccd1 vccd1 _3229_ sky130_fd_sc_hd__buf_2
X_8518_ reg_data\[1\]\[0\] _3118_ _4180_ vssd1 vssd1 vccd1 vccd1 _4181_ sky130_fd_sc_hd__mux2_1
X_9498_ clknet_leaf_11_i_clk _0642_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8449_ _4143_ vssd1 vssd1 vccd1 vccd1 _4144_ sky130_fd_sc_hd__buf_4
X_7820_ _3794_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__clkbuf_1
X_7751_ _3218_ reg_data\[26\]\[8\] _3749_ vssd1 vssd1 vccd1 vccd1 _3758_ sky130_fd_sc_hd__mux2_1
X_4963_ reg_data\[5\]\[8\] _1179_ _1285_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__and3_1
X_6702_ i_data[22] vssd1 vssd1 vccd1 vccd1 _3175_ sky130_fd_sc_hd__clkbuf_4
X_7682_ _3721_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__clkbuf_1
X_6633_ _3125_ _3127_ vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__nor2_4
X_4894_ _1506_ vssd1 vssd1 vccd1 vccd1 rdata1\[7\] sky130_fd_sc_hd__clkbuf_2
X_9421_ clknet_leaf_49_i_clk _0565_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_9352_ clknet_leaf_52_i_clk _0496_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6564_ _3087_ vssd1 vssd1 vccd1 vccd1 o_data2[3] sky130_fd_sc_hd__buf_2
X_8303_ _3917_ reg_data\[15\]\[28\] _4057_ vssd1 vssd1 vccd1 vccd1 _4066_ sky130_fd_sc_hd__mux2_1
X_9283_ clknet_leaf_61_i_clk _0427_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_5515_ reg_data\[1\]\[17\] _1729_ _1793_ _1794_ reg_data\[15\]\[17\] vssd1 vssd1
+ vccd1 vccd1 _2108_ sky130_fd_sc_hd__a32o_1
X_6495_ _3050_ vssd1 vssd1 vccd1 vccd1 o_data1[3] sky130_fd_sc_hd__buf_2
X_8234_ _4029_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__clkbuf_1
X_5446_ reg_data\[0\]\[16\] _1775_ _2038_ _2039_ _2040_ vssd1 vssd1 vccd1 vccd1 _2041_
+ sky130_fd_sc_hd__a2111o_1
X_8165_ _3915_ reg_data\[13\]\[27\] _3985_ vssd1 vssd1 vccd1 vccd1 _3993_ sky130_fd_sc_hd__mux2_1
X_5377_ reg_data\[17\]\[15\] _1766_ _1708_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__and3_1
X_8096_ _3915_ reg_data\[30\]\[27\] _3948_ vssd1 vssd1 vccd1 vccd1 _3956_ sky130_fd_sc_hd__mux2_1
X_7116_ _3125_ _3418_ vssd1 vssd1 vccd1 vccd1 _3419_ sky130_fd_sc_hd__nor2_4
X_7047_ _3381_ _3307_ vssd1 vssd1 vccd1 vccd1 _3382_ sky130_fd_sc_hd__nand2_4
X_8998_ clknet_leaf_48_i_clk _0142_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_7949_ i_data[3] vssd1 vssd1 vccd1 vccd1 _3865_ sky130_fd_sc_hd__clkbuf_4
X_9619_ clknet_leaf_31_i_clk _0763_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5300_ reg_data\[23\]\[13\] _1834_ _1835_ reg_data\[19\]\[13\] vssd1 vssd1 vccd1
+ vccd1 _1900_ sky130_fd_sc_hd__a22o_1
X_6280_ reg_data\[13\]\[30\] _2473_ _1086_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__and3_1
X_5231_ _1198_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__clkbuf_4
X_5162_ reg_data\[22\]\[12\] _1536_ _1651_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__and3_1
X_5093_ reg_data\[2\]\[10\] _1002_ _1295_ _1296_ reg_data\[11\]\[10\] vssd1 vssd1
+ vccd1 vccd1 _1699_ sky130_fd_sc_hd__a32o_1
X_8921_ clknet_leaf_1_i_clk _0065_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8852_ reg_data\[11\]\[30\] i_data[30] _4323_ vssd1 vssd1 vccd1 vccd1 _4357_ sky130_fd_sc_hd__mux2_1
X_8783_ _4320_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__clkbuf_1
X_7803_ _3195_ reg_data\[27\]\[0\] _3785_ vssd1 vssd1 vccd1 vccd1 _3786_ sky130_fd_sc_hd__mux2_1
X_5995_ reg_data\[24\]\[24\] _2453_ _2454_ reg_data\[28\]\[24\] _2572_ vssd1 vssd1
+ vccd1 vccd1 _2573_ sky130_fd_sc_hd__a221o_1
X_7734_ _3748_ vssd1 vssd1 vccd1 vccd1 _3749_ sky130_fd_sc_hd__buf_4
X_4946_ reg_data\[27\]\[8\] _1096_ _1554_ _1555_ _1556_ vssd1 vssd1 vccd1 vccd1 _1557_
+ sky130_fd_sc_hd__a2111o_1
X_7665_ _3601_ _3675_ vssd1 vssd1 vccd1 vccd1 _3712_ sky130_fd_sc_hd__nand2_2
X_4877_ _1067_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__clkbuf_4
X_6616_ _3114_ vssd1 vssd1 vccd1 vccd1 o_data2[28] sky130_fd_sc_hd__buf_2
X_9404_ clknet_leaf_71_i_clk _0548_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_7596_ i_rd[3] i_rd[4] _3119_ _3120_ vssd1 vssd1 vccd1 vccd1 _3675_ sky130_fd_sc_hd__and4_4
X_9335_ clknet_leaf_25_i_clk _0479_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6547_ _3077_ vssd1 vssd1 vccd1 vccd1 o_data1[28] sky130_fd_sc_hd__buf_2
X_9266_ clknet_leaf_35_i_clk _0410_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6478_ reg_data\[27\]\[1\] _1198_ _3035_ _3036_ _3037_ vssd1 vssd1 vccd1 vccd1 _3038_
+ sky130_fd_sc_hd__a2111o_1
X_9197_ clknet_leaf_32_i_clk _0341_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_8217_ _4020_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__clkbuf_1
X_5429_ reg_data\[8\]\[15\] _1841_ _1842_ reg_data\[10\]\[15\] _2024_ vssd1 vssd1
+ vccd1 vccd1 _2025_ sky130_fd_sc_hd__a221o_1
X_8148_ _3898_ reg_data\[13\]\[19\] _3974_ vssd1 vssd1 vccd1 vccd1 _3984_ sky130_fd_sc_hd__mux2_1
X_8079_ _3898_ reg_data\[30\]\[19\] _3937_ vssd1 vssd1 vccd1 vccd1 _3947_ sky130_fd_sc_hd__mux2_1
X_4800_ reg_data\[23\]\[5\] _1206_ _1209_ reg_data\[19\]\[5\] vssd1 vssd1 vccd1 vccd1
+ _1416_ sky130_fd_sc_hd__a22o_1
X_5780_ reg_data\[27\]\[21\] _1833_ _2361_ _2362_ _2363_ vssd1 vssd1 vccd1 vccd1 _2364_
+ sky130_fd_sc_hd__a2111o_1
X_4731_ reg_data\[4\]\[4\] _1177_ _1283_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__and3_1
X_7450_ _3596_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__clkbuf_1
X_4662_ reg_data\[6\]\[3\] _1175_ _1152_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__and3_1
X_6401_ reg_data\[24\]\[0\] _1126_ _1129_ reg_data\[28\]\[0\] _2963_ vssd1 vssd1 vccd1
+ vccd1 _2964_ sky130_fd_sc_hd__a221o_1
X_7381_ reg_data\[3\]\[28\] _3187_ _3551_ vssd1 vssd1 vccd1 vccd1 _3560_ sky130_fd_sc_hd__mux2_1
X_4593_ rs2_mux\[0\] _1006_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__nor2_1
X_9120_ clknet_leaf_2_i_clk _0264_ vssd1 vssd1 vccd1 vccd1 reg_data\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6332_ reg_data\[5\]\[31\] _1085_ _2530_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__and3_1
X_6263_ reg_data\[8\]\[29\] _2447_ _2448_ reg_data\[10\]\[29\] _2830_ vssd1 vssd1
+ vccd1 vccd1 _2831_ sky130_fd_sc_hd__a221o_1
X_9051_ clknet_leaf_4_i_clk _0195_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5214_ _1142_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__buf_2
X_8002_ _3858_ vssd1 vssd1 vccd1 vccd1 _3901_ sky130_fd_sc_hd__buf_4
X_6194_ reg_data\[3\]\[28\] _2421_ _2761_ _2762_ _2763_ vssd1 vssd1 vccd1 vccd1 _2764_
+ sky130_fd_sc_hd__a2111o_1
X_5145_ reg_data\[0\]\[11\] _1174_ _1746_ _1747_ _1748_ vssd1 vssd1 vccd1 vccd1 _1749_
+ sky130_fd_sc_hd__a2111o_1
X_5076_ reg_data\[17\]\[10\] _1509_ _1275_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__and3_1
X_8904_ clknet_leaf_49_i_clk _0048_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_9884_ clknet_leaf_34_i_clk _0954_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_8835_ _4348_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__clkbuf_1
X_5978_ reg_data\[6\]\[24\] _2555_ _2237_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__and3_1
X_8766_ _3903_ reg_data\[29\]\[21\] _4310_ vssd1 vssd1 vccd1 vccd1 _4312_ sky130_fd_sc_hd__mux2_1
X_7717_ _3252_ reg_data\[25\]\[24\] _3735_ vssd1 vssd1 vccd1 vccd1 _3740_ sky130_fd_sc_hd__mux2_1
X_8697_ _4275_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__clkbuf_1
X_4929_ reg_data\[25\]\[8\] _1037_ _1537_ _1538_ _1539_ vssd1 vssd1 vccd1 vccd1 _1540_
+ sky130_fd_sc_hd__a2111o_1
X_7648_ _3703_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__clkbuf_1
X_7579_ _3666_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__clkbuf_1
X_9318_ clknet_leaf_51_i_clk _0462_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_9249_ clknet_leaf_1_i_clk _0393_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6950_ _3241_ reg_data\[10\]\[19\] _3320_ vssd1 vssd1 vccd1 vccd1 _3330_ sky130_fd_sc_hd__mux2_1
X_5901_ reg_data\[27\]\[23\] _2392_ _2479_ _2480_ _2481_ vssd1 vssd1 vccd1 vccd1 _2482_
+ sky130_fd_sc_hd__a2111o_1
X_6881_ _3292_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__clkbuf_1
X_5832_ _2391_ _2402_ _2408_ _2414_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__or4_1
X_8620_ _4234_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__clkbuf_1
X_5763_ reg_data\[25\]\[21\] _1810_ _2344_ _2345_ _2346_ vssd1 vssd1 vccd1 vccd1 _2347_
+ sky130_fd_sc_hd__a2111o_1
X_8551_ reg_data\[1\]\[16\] _3162_ _4191_ vssd1 vssd1 vccd1 vccd1 _4198_ sky130_fd_sc_hd__mux2_1
X_7502_ _3602_ vssd1 vssd1 vccd1 vccd1 _3625_ sky130_fd_sc_hd__buf_4
X_4714_ reg_data\[26\]\[4\] _1132_ _1134_ reg_data\[29\]\[4\] vssd1 vssd1 vccd1 vccd1
+ _1333_ sky130_fd_sc_hd__a22o_1
X_5694_ reg_data\[8\]\[20\] _1797_ _1798_ reg_data\[10\]\[20\] _2280_ vssd1 vssd1
+ vccd1 vccd1 _2281_ sky130_fd_sc_hd__a221o_1
X_8482_ _4161_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__clkbuf_1
X_7433_ _3243_ reg_data\[20\]\[20\] _3587_ vssd1 vssd1 vccd1 vccd1 _3588_ sky130_fd_sc_hd__mux2_1
X_4645_ reg_data\[8\]\[3\] _1116_ _1119_ reg_data\[10\]\[3\] _1265_ vssd1 vssd1 vccd1
+ vccd1 _1266_ sky130_fd_sc_hd__a221o_1
X_7364_ _3528_ vssd1 vssd1 vccd1 vccd1 _3551_ sky130_fd_sc_hd__buf_4
X_4576_ _1166_ _1197_ _1156_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__and3_4
X_9103_ clknet_leaf_30_i_clk _0247_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6315_ reg_data\[27\]\[30\] _2439_ _2878_ _2879_ _2880_ vssd1 vssd1 vccd1 vccd1 _2881_
+ sky130_fd_sc_hd__a2111o_1
X_7295_ _3514_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__clkbuf_1
X_9034_ clknet_leaf_50_i_clk _0178_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6246_ reg_data\[20\]\[29\] _1146_ _1160_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__and3_1
X_6177_ reg_data\[23\]\[28\] _2393_ _2394_ reg_data\[19\]\[28\] vssd1 vssd1 vccd1
+ vccd1 _2748_ sky130_fd_sc_hd__a22o_1
X_5128_ reg_data\[8\]\[11\] _1116_ _1119_ reg_data\[10\]\[11\] _1732_ vssd1 vssd1
+ vccd1 vccd1 _1733_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_54_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5059_ reg_data\[12\]\[10\] _1381_ _1606_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__and3_1
X_9867_ clknet_leaf_72_i_clk _0937_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_69_i_clk clknet_3_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_8818_ _4339_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__clkbuf_1
X_9798_ clknet_leaf_54_i_clk rdata1\[14\] vssd1 vssd1 vccd1 vccd1 r_data1\[14\] sky130_fd_sc_hd__dfxtp_1
X_8749_ _3886_ reg_data\[29\]\[13\] _4299_ vssd1 vssd1 vccd1 vccd1 _4303_ sky130_fd_sc_hd__mux2_1
X_4430_ _1019_ _1051_ _1052_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__and3_1
X_6100_ reg_data\[16\]\[26\] _2449_ _2450_ reg_data\[9\]\[26\] vssd1 vssd1 vccd1 vccd1
+ _2674_ sky130_fd_sc_hd__a22o_1
X_4361_ _0993_ vssd1 vssd1 vccd1 vccd1 rs2_mux\[0\] sky130_fd_sc_hd__clkinv_2
X_7080_ _3233_ reg_data\[8\]\[15\] _3394_ vssd1 vssd1 vccd1 vccd1 _3400_ sky130_fd_sc_hd__mux2_1
X_6031_ reg_data\[20\]\[25\] _2234_ _1283_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__and3_1
X_7982_ _3887_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__clkbuf_1
X_9721_ clknet_leaf_12_i_clk _0865_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6933_ _3321_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__clkbuf_1
X_9652_ clknet_leaf_21_i_clk _0796_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6864_ reg_data\[2\]\[11\] _3152_ _3282_ vssd1 vssd1 vccd1 vccd1 _3284_ sky130_fd_sc_hd__mux2_1
X_5815_ reg_data\[2\]\[22\] _2219_ _2396_ _2397_ reg_data\[11\]\[22\] vssd1 vssd1
+ vccd1 vccd1 _2398_ sky130_fd_sc_hd__a32o_1
X_8603_ _4225_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__clkbuf_1
X_9583_ clknet_leaf_32_i_clk _0727_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6795_ _3239_ reg_data\[22\]\[18\] _3223_ vssd1 vssd1 vccd1 vccd1 _3240_ sky130_fd_sc_hd__mux2_1
X_5746_ reg_data\[13\]\[21\] _2214_ _2102_ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__and3_1
X_8534_ reg_data\[1\]\[8\] _3145_ _4180_ vssd1 vssd1 vccd1 vccd1 _4189_ sky130_fd_sc_hd__mux2_1
X_5677_ reg_data\[20\]\[20\] _2204_ _2035_ vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__and3_1
X_8465_ _4152_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__clkbuf_1
X_4628_ reg_data\[4\]\[3\] _1074_ _1248_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__and3_1
X_7416_ _3227_ reg_data\[20\]\[12\] _3576_ vssd1 vssd1 vccd1 vccd1 _3579_ sky130_fd_sc_hd__mux2_1
X_8396_ _3873_ reg_data\[17\]\[7\] _4108_ vssd1 vssd1 vccd1 vccd1 _4116_ sky130_fd_sc_hd__mux2_1
X_4559_ reg_data\[4\]\[2\] _1179_ _1180_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__and3_1
X_7347_ _3542_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__clkbuf_1
X_7278_ reg_data\[5\]\[11\] _3152_ _3504_ vssd1 vssd1 vccd1 vccd1 _3506_ sky130_fd_sc_hd__mux2_1
X_6229_ reg_data\[7\]\[29\] _2386_ _2795_ _2796_ _2797_ vssd1 vssd1 vccd1 vccd1 _2798_
+ sky130_fd_sc_hd__a2111o_1
X_9017_ clknet_leaf_68_i_clk _0161_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_9919_ clknet_leaf_37_i_clk _0989_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_5600_ reg_data\[2\]\[18\] _1837_ _1901_ _1902_ reg_data\[11\]\[18\] vssd1 vssd1
+ vccd1 vccd1 _2190_ sky130_fd_sc_hd__a32o_1
X_6580_ r_data2\[11\] _3094_ vssd1 vssd1 vccd1 vccd1 _3096_ sky130_fd_sc_hd__and2_1
X_5531_ reg_data\[20\]\[17\] _1629_ _1743_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__and3_1
X_8250_ _4038_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__clkbuf_1
X_7201_ _3464_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_1
X_5462_ reg_data\[22\]\[16\] _1679_ _1622_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__and3_1
X_4413_ _1034_ _1035_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__and2_2
X_8181_ _3863_ reg_data\[14\]\[2\] _3999_ vssd1 vssd1 vccd1 vccd1 _4002_ sky130_fd_sc_hd__mux2_1
X_5393_ _1976_ _1980_ _1984_ _1989_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__or4_1
X_7132_ reg_data\[7\]\[7\] _3143_ _3420_ vssd1 vssd1 vccd1 vccd1 _3428_ sky130_fd_sc_hd__mux2_1
X_7063_ _3216_ reg_data\[8\]\[7\] _3383_ vssd1 vssd1 vccd1 vccd1 _3391_ sky130_fd_sc_hd__mux2_1
X_6014_ _2578_ _2582_ _2586_ _2590_ vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__or4_2
X_9704_ clknet_leaf_56_i_clk _0848_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_7965_ _3875_ reg_data\[9\]\[8\] _3859_ vssd1 vssd1 vccd1 vccd1 _3876_ sky130_fd_sc_hd__mux2_1
X_7896_ _3835_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__clkbuf_1
X_6916_ _3312_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__clkbuf_1
X_6847_ reg_data\[2\]\[3\] _3135_ _3271_ vssd1 vssd1 vccd1 vccd1 _3275_ sky130_fd_sc_hd__mux2_1
X_9635_ clknet_leaf_65_i_clk _0779_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_9566_ clknet_leaf_76_i_clk _0710_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6778_ _3228_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__clkbuf_1
X_5729_ _2314_ vssd1 vssd1 vccd1 vccd1 rdata2\[20\] sky130_fd_sc_hd__clkbuf_1
X_8517_ _4179_ vssd1 vssd1 vccd1 vccd1 _4180_ sky130_fd_sc_hd__buf_4
X_9497_ clknet_leaf_12_i_clk _0641_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8448_ _3200_ _4070_ vssd1 vssd1 vccd1 vccd1 _4143_ sky130_fd_sc_hd__nand2_4
X_8379_ _4106_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__clkbuf_1
X_7750_ _3757_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__clkbuf_1
X_4962_ reg_data\[4\]\[8\] _1460_ _1407_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__and3_1
X_6701_ _3174_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__clkbuf_1
X_4893_ _1497_ _1501_ _1503_ _1505_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__or4_1
X_7681_ _3216_ reg_data\[25\]\[7\] _3713_ vssd1 vssd1 vccd1 vccd1 _3721_ sky130_fd_sc_hd__mux2_1
X_6632_ i_rd[1] _3126_ i_rd[0] vssd1 vssd1 vccd1 vccd1 _3127_ sky130_fd_sc_hd__or3b_4
X_9420_ clknet_leaf_49_i_clk _0564_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_9351_ clknet_leaf_58_i_clk _0495_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6563_ r_data2\[3\] _3083_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__and2_1
X_8302_ _4065_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__clkbuf_1
X_5514_ reg_data\[2\]\[17\] _1613_ _1790_ _1791_ reg_data\[11\]\[17\] vssd1 vssd1
+ vccd1 vccd1 _2107_ sky130_fd_sc_hd__a32o_1
X_6494_ r_data1\[3\] _3046_ vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__and2_1
X_9282_ clknet_leaf_62_i_clk _0426_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8233_ _3915_ reg_data\[14\]\[27\] _4021_ vssd1 vssd1 vccd1 vccd1 _4029_ sky130_fd_sc_hd__mux2_1
X_5445_ reg_data\[5\]\[16\] _1490_ _1925_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__and3_1
X_8164_ _3992_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__clkbuf_1
X_7115_ i_rd[0] i_rd[1] _3126_ vssd1 vssd1 vccd1 vccd1 _3418_ sky130_fd_sc_hd__or3_2
X_5376_ reg_data\[22\]\[15\] _1536_ _1651_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__and3_1
X_8095_ _3955_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__clkbuf_1
X_7046_ _3380_ vssd1 vssd1 vccd1 vccd1 _3381_ sky130_fd_sc_hd__clkbuf_4
X_8997_ clknet_leaf_63_i_clk _0141_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_7948_ _3864_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__clkbuf_1
X_9618_ clknet_leaf_31_i_clk _0762_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_7879_ _3826_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__clkbuf_1
X_9549_ clknet_leaf_16_i_clk _0693_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5230_ _1814_ _1820_ _1826_ _1831_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__or4_1
X_5161_ _1036_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__buf_4
X_5092_ reg_data\[23\]\[10\] _1206_ _1209_ reg_data\[19\]\[10\] vssd1 vssd1 vccd1
+ vccd1 _1698_ sky130_fd_sc_hd__a22o_1
X_8920_ clknet_leaf_62_i_clk _0064_ vssd1 vssd1 vccd1 vccd1 reg_data\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8851_ _4356_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__clkbuf_1
X_5994_ reg_data\[26\]\[24\] _2455_ _2456_ reg_data\[29\]\[24\] vssd1 vssd1 vccd1
+ vccd1 _2572_ sky130_fd_sc_hd__a22o_1
X_8782_ _3919_ reg_data\[29\]\[29\] _4310_ vssd1 vssd1 vccd1 vccd1 _4320_ sky130_fd_sc_hd__mux2_1
X_7802_ _3784_ vssd1 vssd1 vccd1 vccd1 _3785_ sky130_fd_sc_hd__buf_4
X_7733_ _3200_ _3675_ vssd1 vssd1 vccd1 vccd1 _3748_ sky130_fd_sc_hd__nand2_4
X_4945_ reg_data\[1\]\[8\] _1022_ _1109_ _1111_ reg_data\[15\]\[8\] vssd1 vssd1 vccd1
+ vccd1 _1556_ sky130_fd_sc_hd__a32o_1
X_7664_ _3711_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__clkbuf_1
X_4876_ reg_data\[5\]\[7\] _1074_ _1044_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__and3_1
X_6615_ r_data2\[28\] _3105_ vssd1 vssd1 vccd1 vccd1 _3114_ sky130_fd_sc_hd__and2_1
X_7595_ _3674_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__clkbuf_1
X_9403_ clknet_leaf_71_i_clk _0547_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_9334_ clknet_leaf_23_i_clk _0478_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6546_ r_data1\[28\] _3068_ vssd1 vssd1 vccd1 vccd1 _3077_ sky130_fd_sc_hd__and2_1
X_9265_ clknet_leaf_36_i_clk _0409_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6477_ reg_data\[1\]\[1\] _1202_ _1203_ reg_data\[15\]\[1\] vssd1 vssd1 vccd1 vccd1
+ _3037_ sky130_fd_sc_hd__a22o_1
X_9196_ clknet_leaf_28_i_clk _0340_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8216_ _3898_ reg_data\[14\]\[19\] _4010_ vssd1 vssd1 vccd1 vccd1 _4020_ sky130_fd_sc_hd__mux2_1
X_5428_ reg_data\[16\]\[15\] _1843_ _1844_ reg_data\[9\]\[15\] vssd1 vssd1 vccd1 vccd1
+ _2024_ sky130_fd_sc_hd__a22o_1
X_8147_ _3983_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__clkbuf_1
X_5359_ reg_data\[13\]\[14\] _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__and3_1
X_8078_ _3946_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__clkbuf_1
X_7029_ reg_data\[0\]\[24\] _3179_ _3367_ vssd1 vssd1 vccd1 vccd1 _3372_ sky130_fd_sc_hd__mux2_1
X_4730_ reg_data\[6\]\[4\] _1347_ _1152_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__and3_1
X_4661_ reg_data\[3\]\[3\] _1158_ _1278_ _1279_ _1280_ vssd1 vssd1 vccd1 vccd1 _1281_
+ sky130_fd_sc_hd__a2111o_1
X_7380_ _3559_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__clkbuf_1
X_6400_ reg_data\[26\]\[0\] _1131_ _1133_ reg_data\[29\]\[0\] vssd1 vssd1 vccd1 vccd1
+ _2963_ sky130_fd_sc_hd__a22o_1
X_6331_ reg_data\[4\]\[31\] _1072_ _2469_ vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__and3_1
X_4592_ _1213_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__clkbuf_4
X_6262_ reg_data\[16\]\[29\] _2449_ _2450_ reg_data\[9\]\[29\] vssd1 vssd1 vccd1 vccd1
+ _2830_ sky130_fd_sc_hd__a22o_1
X_9050_ clknet_leaf_12_i_clk _0194_ vssd1 vssd1 vccd1 vccd1 reg_data\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6193_ reg_data\[30\]\[28\] _2234_ _1164_ vssd1 vssd1 vccd1 vccd1 _2763_ sky130_fd_sc_hd__and3_1
X_5213_ _1157_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__clkbuf_4
X_8001_ i_data[20] vssd1 vssd1 vccd1 vccd1 _3900_ sky130_fd_sc_hd__clkbuf_4
X_5144_ reg_data\[5\]\[11\] _1179_ _1285_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__and3_1
X_5075_ reg_data\[21\]\[10\] _1272_ _1273_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__and3_1
X_9883_ clknet_leaf_34_i_clk _0953_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_8903_ clknet_leaf_48_i_clk _0047_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8834_ reg_data\[11\]\[21\] i_data[21] _4346_ vssd1 vssd1 vccd1 vccd1 _4348_ sky130_fd_sc_hd__mux2_1
X_5977_ _0999_ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__buf_2
X_8765_ _4311_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__clkbuf_1
X_7716_ _3739_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__clkbuf_1
X_8696_ reg_data\[19\]\[20\] _3170_ _4274_ vssd1 vssd1 vccd1 vccd1 _4275_ sky130_fd_sc_hd__mux2_1
X_4928_ reg_data\[21\]\[8\] _1480_ _1240_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__and3_1
X_7647_ _3250_ reg_data\[24\]\[23\] _3699_ vssd1 vssd1 vccd1 vccd1 _3703_ sky130_fd_sc_hd__mux2_1
X_4859_ reg_data\[16\]\[6\] _1219_ _1221_ reg_data\[9\]\[6\] vssd1 vssd1 vccd1 vccd1
+ _1473_ sky130_fd_sc_hd__a22o_1
X_7578_ reg_data\[23\]\[23\] _3177_ _3662_ vssd1 vssd1 vccd1 vccd1 _3666_ sky130_fd_sc_hd__mux2_1
X_9317_ clknet_leaf_63_i_clk _0461_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6529_ _3045_ vssd1 vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__dlymetal6s2s_1
X_9248_ clknet_leaf_75_i_clk _0392_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_9179_ clknet_leaf_1_i_clk _0323_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5900_ reg_data\[1\]\[23\] _2336_ _2399_ _2400_ reg_data\[15\]\[23\] vssd1 vssd1
+ vccd1 vccd1 _2481_ sky130_fd_sc_hd__a32o_1
X_6880_ reg_data\[2\]\[19\] _3168_ _3282_ vssd1 vssd1 vccd1 vccd1 _3292_ sky130_fd_sc_hd__mux2_1
X_5831_ reg_data\[24\]\[22\] _2409_ _2410_ reg_data\[28\]\[22\] _2413_ vssd1 vssd1
+ vccd1 vccd1 _2414_ sky130_fd_sc_hd__a221o_1
X_5762_ reg_data\[21\]\[21\] _2117_ _1510_ vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__and3_1
X_8550_ _4197_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__clkbuf_1
X_4713_ reg_data\[8\]\[4\] _1116_ _1119_ reg_data\[10\]\[4\] _1331_ vssd1 vssd1 vccd1
+ vccd1 _1332_ sky130_fd_sc_hd__a221o_1
X_7501_ _3624_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__clkbuf_1
X_5693_ reg_data\[16\]\[20\] _1799_ _1800_ reg_data\[9\]\[20\] vssd1 vssd1 vccd1 vccd1
+ _2280_ sky130_fd_sc_hd__a22o_1
X_8481_ _3890_ reg_data\[18\]\[15\] _4155_ vssd1 vssd1 vccd1 vccd1 _4161_ sky130_fd_sc_hd__mux2_1
X_7432_ _3564_ vssd1 vssd1 vccd1 vccd1 _3587_ sky130_fd_sc_hd__buf_4
X_4644_ reg_data\[16\]\[3\] _1121_ _1123_ reg_data\[9\]\[3\] vssd1 vssd1 vccd1 vccd1
+ _1265_ sky130_fd_sc_hd__a22o_1
X_4575_ rs2_mux\[2\] _1013_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__nor2_2
X_7363_ _3550_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__clkbuf_1
X_9102_ clknet_leaf_29_i_clk _0246_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_7294_ reg_data\[5\]\[19\] _3168_ _3504_ vssd1 vssd1 vccd1 vccd1 _3514_ sky130_fd_sc_hd__mux2_1
X_6314_ reg_data\[1\]\[30\] _2510_ _2511_ reg_data\[15\]\[30\] vssd1 vssd1 vccd1 vccd1
+ _2880_ sky130_fd_sc_hd__a22o_1
X_6245_ reg_data\[18\]\[29\] _2422_ _1167_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__and3_1
X_9033_ clknet_leaf_52_i_clk _0177_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6176_ _2734_ _2738_ _2742_ _2746_ vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__or4_2
X_5127_ reg_data\[16\]\[11\] _1121_ _1123_ reg_data\[9\]\[11\] vssd1 vssd1 vccd1 vccd1
+ _1732_ sky130_fd_sc_hd__a22o_1
X_5058_ reg_data\[14\]\[10\] _1253_ _1379_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__and3_1
X_9866_ clknet_leaf_70_i_clk _0936_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8817_ reg_data\[11\]\[13\] i_data[13] _4335_ vssd1 vssd1 vccd1 vccd1 _4339_ sky130_fd_sc_hd__mux2_1
X_9797_ clknet_leaf_54_i_clk rdata1\[13\] vssd1 vssd1 vccd1 vccd1 r_data1\[13\] sky130_fd_sc_hd__dfxtp_1
X_8748_ _4302_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__clkbuf_1
X_8679_ reg_data\[19\]\[12\] _3154_ _4263_ vssd1 vssd1 vccd1 vccd1 _4266_ sky130_fd_sc_hd__mux2_1
X_4360_ _0992_ i_rs2[0] i_rs_valid vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__mux2_2
X_6030_ reg_data\[30\]\[25\] _1146_ _2006_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__and3_1
X_7981_ _3886_ reg_data\[9\]\[13\] _3880_ vssd1 vssd1 vccd1 vccd1 _3887_ sky130_fd_sc_hd__mux2_1
X_9720_ clknet_leaf_13_i_clk _0864_ vssd1 vssd1 vccd1 vccd1 reg_data\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6932_ _3222_ reg_data\[10\]\[10\] _3320_ vssd1 vssd1 vccd1 vccd1 _3321_ sky130_fd_sc_hd__mux2_1
X_9651_ clknet_leaf_21_i_clk _0795_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6863_ _3283_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__clkbuf_1
X_5814_ _1105_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__clkbuf_4
X_8602_ _3875_ reg_data\[12\]\[8\] _4216_ vssd1 vssd1 vccd1 vccd1 _4225_ sky130_fd_sc_hd__mux2_1
X_9582_ clknet_leaf_39_i_clk _0726_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6794_ i_data[18] vssd1 vssd1 vccd1 vccd1 _3239_ sky130_fd_sc_hd__clkbuf_4
X_5745_ reg_data\[12\]\[21\] _1986_ _2271_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__and3_1
X_8533_ _4188_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__clkbuf_1
X_5676_ reg_data\[30\]\[20\] _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__and3_1
X_8464_ _3873_ reg_data\[18\]\[7\] _4144_ vssd1 vssd1 vccd1 vccd1 _4152_ sky130_fd_sc_hd__mux2_1
X_4627_ _1059_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__clkbuf_4
X_7415_ _3578_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__clkbuf_1
X_8395_ _4115_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__clkbuf_1
X_4558_ _1160_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__buf_4
X_7346_ reg_data\[3\]\[11\] _3152_ _3540_ vssd1 vssd1 vccd1 vccd1 _3542_ sky130_fd_sc_hd__mux2_1
X_4489_ reg_data\[1\]\[2\] _1022_ _1109_ _1111_ reg_data\[15\]\[2\] vssd1 vssd1 vccd1
+ vccd1 _1112_ sky130_fd_sc_hd__a32o_1
X_7277_ _3505_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__clkbuf_1
X_6228_ reg_data\[13\]\[29\] _1076_ _1087_ vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__and3_1
X_9016_ clknet_leaf_69_i_clk _0160_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6159_ _2730_ vssd1 vssd1 vccd1 vccd1 rdata2\[27\] sky130_fd_sc_hd__clkbuf_1
X_9918_ clknet_leaf_32_i_clk _0988_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_9849_ clknet_leaf_24_i_clk rs1_mux\[1\] vssd1 vssd1 vccd1 vccd1 rs1\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_53_i_clk clknet_3_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5530_ reg_data\[30\]\[17\] _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__and3_1
X_5461_ _2055_ vssd1 vssd1 vccd1 vccd1 rdata1\[16\] sky130_fd_sc_hd__clkbuf_1
X_4412_ rs1_mux\[0\] _1026_ _1030_ rs1_mux\[3\] vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__and4_1
X_7200_ reg_data\[6\]\[7\] _3143_ _3456_ vssd1 vssd1 vccd1 vccd1 _3464_ sky130_fd_sc_hd__mux2_1
X_8180_ _4001_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__clkbuf_1
X_5392_ reg_data\[7\]\[15\] _1780_ _1985_ _1987_ _1988_ vssd1 vssd1 vccd1 vccd1 _1989_
+ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_68_i_clk clknet_3_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_7131_ _3427_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_1
X_7062_ _3390_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_1
X_6013_ reg_data\[7\]\[25\] _2386_ _2587_ _2588_ _2589_ vssd1 vssd1 vccd1 vccd1 _2590_
+ sky130_fd_sc_hd__a2111o_1
X_7964_ i_data[8] vssd1 vssd1 vccd1 vccd1 _3875_ sky130_fd_sc_hd__clkbuf_4
X_9703_ clknet_leaf_56_i_clk _0847_ vssd1 vssd1 vccd1 vccd1 reg_data\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6915_ _3206_ reg_data\[10\]\[2\] _3309_ vssd1 vssd1 vccd1 vccd1 _3312_ sky130_fd_sc_hd__mux2_1
X_7895_ _3225_ reg_data\[28\]\[11\] _3833_ vssd1 vssd1 vccd1 vccd1 _3835_ sky130_fd_sc_hd__mux2_1
X_6846_ _3274_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__clkbuf_1
X_9634_ clknet_leaf_65_i_clk _0778_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_9565_ clknet_leaf_0_i_clk _0709_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6777_ _3227_ reg_data\[22\]\[12\] _3223_ vssd1 vssd1 vccd1 vccd1 _3228_ sky130_fd_sc_hd__mux2_1
X_8516_ _3269_ _3491_ vssd1 vssd1 vccd1 vccd1 _4179_ sky130_fd_sc_hd__nor2_4
X_5728_ _2305_ _2309_ _2311_ _2313_ vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__or4_1
X_9496_ clknet_leaf_13_i_clk _0640_ vssd1 vssd1 vccd1 vccd1 reg_data\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8447_ _4142_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__clkbuf_1
X_5659_ reg_data\[23\]\[19\] _1834_ _1835_ reg_data\[19\]\[19\] vssd1 vssd1 vccd1
+ vccd1 _2247_ sky130_fd_sc_hd__a22o_1
X_8378_ _3923_ reg_data\[16\]\[31\] _4071_ vssd1 vssd1 vccd1 vccd1 _4106_ sky130_fd_sc_hd__mux2_1
X_7329_ reg_data\[3\]\[3\] _3135_ _3529_ vssd1 vssd1 vccd1 vccd1 _3533_ sky130_fd_sc_hd__mux2_1
X_4961_ reg_data\[6\]\[8\] _1347_ _1152_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__and3_1
X_6700_ reg_data\[4\]\[21\] _3173_ _3171_ vssd1 vssd1 vccd1 vccd1 _3174_ sky130_fd_sc_hd__mux2_1
X_4892_ reg_data\[24\]\[7\] _1127_ _1130_ reg_data\[28\]\[7\] _1504_ vssd1 vssd1 vccd1
+ vccd1 _1505_ sky130_fd_sc_hd__a221o_1
X_7680_ _3720_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__clkbuf_1
X_6631_ i_write i_reset_n vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__nand2_1
X_9350_ clknet_leaf_54_i_clk _0494_ vssd1 vssd1 vccd1 vccd1 reg_data\[26\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8301_ _3915_ reg_data\[15\]\[27\] _4057_ vssd1 vssd1 vccd1 vccd1 _4065_ sky130_fd_sc_hd__mux2_1
X_6562_ _3086_ vssd1 vssd1 vccd1 vccd1 o_data2[2] sky130_fd_sc_hd__buf_2
X_6493_ _3049_ vssd1 vssd1 vccd1 vccd1 o_data1[2] sky130_fd_sc_hd__buf_2
X_5513_ reg_data\[23\]\[17\] _1787_ _1788_ reg_data\[19\]\[17\] vssd1 vssd1 vccd1
+ vccd1 _2106_ sky130_fd_sc_hd__a22o_1
X_9281_ clknet_leaf_67_i_clk _0425_ vssd1 vssd1 vccd1 vccd1 reg_data\[24\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_8232_ _4028_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__clkbuf_1
X_5444_ reg_data\[4\]\[16\] _1718_ _1863_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__and3_1
X_8163_ _3913_ reg_data\[13\]\[26\] _3985_ vssd1 vssd1 vccd1 vccd1 _3992_ sky130_fd_sc_hd__mux2_1
X_7114_ _3417_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
X_5375_ _1972_ vssd1 vssd1 vccd1 vccd1 rdata2\[14\] sky130_fd_sc_hd__clkbuf_1
X_8094_ _3913_ reg_data\[30\]\[26\] _3948_ vssd1 vssd1 vccd1 vccd1 _3955_ sky130_fd_sc_hd__mux2_1
X_7045_ i_rd[1] i_write i_reset_n i_rd[0] vssd1 vssd1 vccd1 vccd1 _3380_ sky130_fd_sc_hd__and4b_1
X_8996_ clknet_leaf_63_i_clk _0140_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_7947_ _3863_ reg_data\[9\]\[2\] _3859_ vssd1 vssd1 vccd1 vccd1 _3864_ sky130_fd_sc_hd__mux2_1
X_7878_ _3208_ reg_data\[28\]\[3\] _3822_ vssd1 vssd1 vccd1 vccd1 _3826_ sky130_fd_sc_hd__mux2_1
X_6829_ _3262_ reg_data\[22\]\[29\] _3244_ vssd1 vssd1 vccd1 vccd1 _3263_ sky130_fd_sc_hd__mux2_1
X_9617_ clknet_leaf_31_i_clk _0761_ vssd1 vssd1 vccd1 vccd1 reg_data\[16\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_9548_ clknet_leaf_23_i_clk _0692_ vssd1 vssd1 vccd1 vccd1 reg_data\[14\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_9479_ clknet_leaf_46_i_clk _0623_ vssd1 vssd1 vccd1 vccd1 reg_data\[30\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_5160_ _1763_ vssd1 vssd1 vccd1 vccd1 rdata2\[11\] sky130_fd_sc_hd__clkbuf_1
X_5091_ _1683_ _1687_ _1691_ _1696_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__or4_1
X_8850_ reg_data\[11\]\[29\] i_data[29] _4346_ vssd1 vssd1 vccd1 vccd1 _4356_ sky130_fd_sc_hd__mux2_1
X_8781_ _4319_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__clkbuf_1
X_5993_ reg_data\[8\]\[24\] _2447_ _2448_ reg_data\[10\]\[24\] _2570_ vssd1 vssd1
+ vccd1 vccd1 _2571_ sky130_fd_sc_hd__a221o_1
X_7801_ _3638_ _3675_ vssd1 vssd1 vccd1 vccd1 _3784_ sky130_fd_sc_hd__nand2_4
X_7732_ _3747_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__clkbuf_1
X_4944_ reg_data\[2\]\[8\] _1103_ _1104_ _1106_ reg_data\[11\]\[8\] vssd1 vssd1 vccd1
+ vccd1 _1555_ sky130_fd_sc_hd__a32o_1
X_7663_ _3266_ reg_data\[24\]\[31\] _3676_ vssd1 vssd1 vccd1 vccd1 _3711_ sky130_fd_sc_hd__mux2_1
X_9402_ clknet_leaf_61_i_clk _0546_ vssd1 vssd1 vccd1 vccd1 reg_data\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_4875_ reg_data\[6\]\[7\] _1072_ _1048_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__and3_1
X_6614_ _3113_ vssd1 vssd1 vccd1 vccd1 o_data2[27] sky130_fd_sc_hd__buf_2
X_7594_ reg_data\[23\]\[31\] _3193_ _3639_ vssd1 vssd1 vccd1 vccd1 _3674_ sky130_fd_sc_hd__mux2_1
X_9333_ clknet_leaf_21_i_clk _0477_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_6__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_6545_ _3076_ vssd1 vssd1 vccd1 vccd1 o_data1[27] sky130_fd_sc_hd__buf_2
X_9264_ clknet_leaf_35_i_clk _0408_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_8215_ _4019_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__clkbuf_1
X_6476_ reg_data\[2\]\[1\] _1001_ _1168_ _1200_ reg_data\[11\]\[1\] vssd1 vssd1 vccd1
+ vccd1 _3036_ sky130_fd_sc_hd__a32o_1
X_9195_ clknet_leaf_44_i_clk _0339_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5427_ reg_data\[27\]\[15\] _1833_ _2020_ _2021_ _2022_ vssd1 vssd1 vccd1 vccd1 _2023_
+ sky130_fd_sc_hd__a2111o_1
X_8146_ _3896_ reg_data\[13\]\[18\] _3974_ vssd1 vssd1 vccd1 vccd1 _3983_ sky130_fd_sc_hd__mux2_1
X_5358_ reg_data\[0\]\[14\] _1821_ _1952_ _1953_ _1955_ vssd1 vssd1 vccd1 vccd1 _1956_
+ sky130_fd_sc_hd__a2111o_1
X_8077_ _3896_ reg_data\[30\]\[18\] _3937_ vssd1 vssd1 vccd1 vccd1 _3946_ sky130_fd_sc_hd__mux2_1
X_7028_ _3371_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__clkbuf_1
X_5289_ reg_data\[20\]\[13\] _1629_ _1743_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__and3_1
X_8979_ clknet_leaf_33_i_clk _0123_ vssd1 vssd1 vccd1 vccd1 reg_data\[10\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_4660_ reg_data\[20\]\[3\] _1166_ _1180_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__and3_1
X_6330_ reg_data\[6\]\[31\] _1020_ _1236_ vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__and3_1
X_4591_ _1001_ _1197_ _1212_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__and3_4
X_6261_ reg_data\[27\]\[29\] _2439_ _2826_ _2827_ _2828_ vssd1 vssd1 vccd1 vccd1 _2829_
+ sky130_fd_sc_hd__a2111o_1
X_6192_ reg_data\[20\]\[28\] _1146_ _1160_ vssd1 vssd1 vccd1 vccd1 _2762_ sky130_fd_sc_hd__and3_1
X_8000_ _3899_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__clkbuf_1
X_5212_ reg_data\[25\]\[12\] _1810_ _1811_ _1812_ _1813_ vssd1 vssd1 vccd1 vccd1 _1814_
+ sky130_fd_sc_hd__a2111o_1
X_5143_ reg_data\[4\]\[11\] _1460_ _1407_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__and3_1
X_5074_ reg_data\[22\]\[10\] _1679_ _1622_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__and3_1
X_9882_ clknet_leaf_31_i_clk _0952_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_8902_ clknet_leaf_51_i_clk _0046_ vssd1 vssd1 vccd1 vccd1 reg_data\[22\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8833_ _4347_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__clkbuf_1
X_5976_ reg_data\[3\]\[24\] _2421_ _2551_ _2552_ _2553_ vssd1 vssd1 vccd1 vccd1 _2554_
+ sky130_fd_sc_hd__a2111o_1
X_8764_ _3900_ reg_data\[29\]\[20\] _4310_ vssd1 vssd1 vccd1 vccd1 _4311_ sky130_fd_sc_hd__mux2_1
X_7715_ _3250_ reg_data\[25\]\[23\] _3735_ vssd1 vssd1 vccd1 vccd1 _3739_ sky130_fd_sc_hd__mux2_1
X_8695_ _4251_ vssd1 vssd1 vccd1 vccd1 _4274_ sky130_fd_sc_hd__buf_4
X_4927_ reg_data\[17\]\[8\] _1042_ _1238_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__and3_1
X_7646_ _3702_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__clkbuf_1
X_4858_ reg_data\[27\]\[6\] _1199_ _1469_ _1470_ _1471_ vssd1 vssd1 vccd1 vccd1 _1472_
+ sky130_fd_sc_hd__a2111o_1
X_7577_ _3665_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__clkbuf_1
X_9316_ clknet_leaf_47_i_clk _0460_ vssd1 vssd1 vccd1 vccd1 reg_data\[25\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_4789_ reg_data\[3\]\[5\] _1158_ _1400_ _1403_ _1404_ vssd1 vssd1 vccd1 vccd1 _1405_
+ sky130_fd_sc_hd__a2111o_1
X_6528_ _3067_ vssd1 vssd1 vccd1 vccd1 o_data1[19] sky130_fd_sc_hd__buf_2
X_6459_ reg_data\[21\]\[1\] _2489_ _1144_ vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__and3_1
X_9247_ clknet_leaf_77_i_clk _0391_ vssd1 vssd1 vccd1 vccd1 reg_data\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_9178_ clknet_leaf_5_i_clk _0322_ vssd1 vssd1 vccd1 vccd1 reg_data\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8129_ _3962_ vssd1 vssd1 vccd1 vccd1 _3974_ sky130_fd_sc_hd__buf_4
X_5830_ reg_data\[26\]\[22\] _2411_ _2412_ reg_data\[29\]\[22\] vssd1 vssd1 vccd1
+ vccd1 _2413_ sky130_fd_sc_hd__a22o_1
X_5761_ reg_data\[17\]\[21\] _1883_ _1395_ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__and3_1
X_4712_ reg_data\[16\]\[4\] _1121_ _1123_ reg_data\[9\]\[4\] vssd1 vssd1 vccd1 vccd1
+ _1331_ sky130_fd_sc_hd__a22o_1
X_8480_ _4160_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__clkbuf_1
X_7500_ _3241_ reg_data\[21\]\[19\] _3614_ vssd1 vssd1 vccd1 vccd1 _3624_ sky130_fd_sc_hd__mux2_1
X_7431_ _3586_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__clkbuf_1
X_5692_ reg_data\[27\]\[20\] _1786_ _2276_ _2277_ _2278_ vssd1 vssd1 vccd1 vccd1 _2279_
+ sky130_fd_sc_hd__a2111o_1
X_4643_ reg_data\[27\]\[3\] _1096_ _1261_ _1262_ _1263_ vssd1 vssd1 vccd1 vccd1 _1264_
+ sky130_fd_sc_hd__a2111o_1
X_7362_ reg_data\[3\]\[19\] _3168_ _3540_ vssd1 vssd1 vccd1 vccd1 _3550_ sky130_fd_sc_hd__mux2_1
X_4574_ _1154_ _1170_ _1182_ _1195_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__or4_2
X_9101_ clknet_leaf_27_i_clk _0245_ vssd1 vssd1 vccd1 vccd1 reg_data\[6\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6313_ reg_data\[2\]\[30\] _2443_ _2507_ _2508_ reg_data\[11\]\[30\] vssd1 vssd1
+ vccd1 vccd1 _2879_ sky130_fd_sc_hd__a32o_1
X_7293_ _3513_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__clkbuf_1
X_6244_ reg_data\[25\]\[29\] _2416_ _2809_ _2810_ _2811_ vssd1 vssd1 vccd1 vccd1 _2812_
+ sky130_fd_sc_hd__a2111o_1
X_9032_ clknet_leaf_53_i_clk _0176_ vssd1 vssd1 vccd1 vccd1 reg_data\[8\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6175_ reg_data\[7\]\[28\] _2386_ _2743_ _2744_ _2745_ vssd1 vssd1 vccd1 vccd1 _2746_
+ sky130_fd_sc_hd__a2111o_1
X_5126_ reg_data\[27\]\[11\] _1096_ _1727_ _1728_ _1730_ vssd1 vssd1 vccd1 vccd1 _1731_
+ sky130_fd_sc_hd__a2111o_1
X_5057_ reg_data\[0\]\[10\] _1070_ _1661_ _1662_ _1663_ vssd1 vssd1 vccd1 vccd1 _1664_
+ sky130_fd_sc_hd__a2111o_1
X_9865_ clknet_leaf_72_i_clk _0935_ vssd1 vssd1 vccd1 vccd1 reg_data\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8816_ _4338_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__clkbuf_1
X_9796_ clknet_leaf_54_i_clk rdata1\[12\] vssd1 vssd1 vccd1 vccd1 r_data1\[12\] sky130_fd_sc_hd__dfxtp_1
X_5959_ reg_data\[23\]\[24\] _2393_ _2394_ reg_data\[19\]\[24\] vssd1 vssd1 vccd1
+ vccd1 _2538_ sky130_fd_sc_hd__a22o_1
X_8747_ _3884_ reg_data\[29\]\[12\] _4299_ vssd1 vssd1 vccd1 vccd1 _4302_ sky130_fd_sc_hd__mux2_1
X_8678_ _4265_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__clkbuf_1
X_7629_ _3693_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__clkbuf_1
X_7980_ i_data[13] vssd1 vssd1 vccd1 vccd1 _3886_ sky130_fd_sc_hd__clkbuf_4
X_6931_ _3308_ vssd1 vssd1 vccd1 vccd1 _3320_ sky130_fd_sc_hd__buf_4
X_9650_ clknet_leaf_30_i_clk _0794_ vssd1 vssd1 vccd1 vccd1 reg_data\[17\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6862_ reg_data\[2\]\[10\] _3149_ _3282_ vssd1 vssd1 vccd1 vccd1 _3283_ sky130_fd_sc_hd__mux2_1
X_9581_ clknet_leaf_40_i_clk _0725_ vssd1 vssd1 vccd1 vccd1 reg_data\[15\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5813_ _1064_ vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__clkbuf_4
X_8601_ _4224_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__clkbuf_1
X_8532_ reg_data\[1\]\[7\] _3143_ _4180_ vssd1 vssd1 vccd1 vccd1 _4188_ sky130_fd_sc_hd__mux2_1
X_6793_ _3238_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__clkbuf_1
X_5744_ reg_data\[14\]\[21\] _1867_ _2156_ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__and3_1
X_5675_ reg_data\[18\]\[20\] _2261_ _2090_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__and3_1
X_8463_ _4151_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__clkbuf_1
X_4626_ reg_data\[6\]\[3\] _1072_ _1048_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__and3_1
X_7414_ _3225_ reg_data\[20\]\[11\] _3576_ vssd1 vssd1 vccd1 vccd1 _3578_ sky130_fd_sc_hd__mux2_1
X_8394_ _3871_ reg_data\[17\]\[6\] _4108_ vssd1 vssd1 vccd1 vccd1 _4115_ sky130_fd_sc_hd__mux2_1
X_7345_ _3541_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__clkbuf_1
X_4557_ _1000_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__clkbuf_4
X_4488_ _1110_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__buf_4
X_7276_ reg_data\[5\]\[10\] _3149_ _3504_ vssd1 vssd1 vccd1 vccd1 _3505_ sky130_fd_sc_hd__mux2_1
X_6227_ reg_data\[12\]\[29\] _1082_ _2271_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__and3_1
X_9015_ clknet_leaf_14_i_clk _0159_ vssd1 vssd1 vccd1 vccd1 reg_data\[0\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6158_ _2721_ _2725_ _2727_ _2729_ vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__or4_1
X_5109_ reg_data\[20\]\[11\] _1597_ _1315_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__and3_1
X_6089_ reg_data\[4\]\[26\] _2430_ _1180_ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__and3_1
X_9917_ clknet_leaf_37_i_clk _0987_ vssd1 vssd1 vccd1 vccd1 reg_data\[11\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_9848_ clknet_leaf_24_i_clk rs1_mux\[0\] vssd1 vssd1 vccd1 vccd1 rs1\[0\] sky130_fd_sc_hd__dfxtp_1
X_9779_ clknet_leaf_35_i_clk _0923_ vssd1 vssd1 vccd1 vccd1 reg_data\[19\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5460_ _2046_ _2050_ _2052_ _2054_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__or4_1
X_4411_ _1017_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__buf_2
X_5391_ reg_data\[12\]\[15\] _1608_ _1128_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__and3_1
X_7130_ reg_data\[7\]\[6\] _3141_ _3420_ vssd1 vssd1 vccd1 vccd1 _3427_ sky130_fd_sc_hd__mux2_1
X_7061_ _3214_ reg_data\[8\]\[6\] _3383_ vssd1 vssd1 vccd1 vccd1 _3390_ sky130_fd_sc_hd__mux2_1
X_6012_ reg_data\[13\]\[25\] _2214_ _2102_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__and3_1
.ends

