
.include ../../elements/inc_lib.spice
.include simulation/rom_dec.spice

.param VCC=1.8

VVCC VCC 0 PWL 0ns 0 1ns 0 1.1ns {VCC}
VVSS VSS 0 PWL 0n 0

.include simulation/stimuli_rom_dec.cir
.options timeint reltol=1e-3 abstol=1e-5
.options linsol type=belos AZ_tol=1.0e-3
.tran 1p 1025n
.print tran format=raw file=simulation/rom_dec.spice.raw v(*)

.GLOBAL VCC
.GLOBAL VSS
.end
