* NGSPICE file created from rv_alu2.ext - technology: sky130A


X_3155_ _0461_ u_bits.i_op2\[26\] _0465_ u_bits.i_op1\[26\] VSS VSS VCC VCC
+ _0959_ sky130_fd_sc_hs__a22o_1
X_3086_ _0849_ _0850_ VSS VSS VCC VCC _0894_ sky130_fd_sc_hs__nand2_1
X_3988_ _1376_ _0909_ _1639_ VSS VSS VCC VCC _1648_ sky130_fd_sc_hs__mux2_1
X_5727_ clknet_leaf_19_i_clk _0370_ VSS VSS VCC VCC u_muldiv.dividend\[11\]
+ sky130_fd_sc_hs__dfxtp_1
X_2939_ u_bits.i_op1\[21\] u_bits.i_op1\[22\] _0657_ VSS VSS VCC VCC _0752_
+ sky130_fd_sc_hs__mux2_1
X_5658_ clknet_leaf_25_i_clk _0301_ VSS VSS VCC VCC u_muldiv.o_div\[4\] sky130_fd_sc_hs__dfxtp_1
X_4609_ u_muldiv.divisor\[21\] u_muldiv.dividend\[21\] VSS VSS VCC VCC _2032_
+ sky130_fd_sc_hs__or2b_1
X_5589_ clknet_leaf_23_i_clk _0236_ VSS VSS VCC VCC u_muldiv.mul\[6\] sky130_fd_sc_hs__dfxtp_1
X_4960_ _2061_ _2065_ _2318_ VSS VSS VCC VCC _2319_ sky130_fd_sc_hs__a21oi_1
X_4891_ u_muldiv.quotient_msk\[3\] _1210_ _2279_ u_muldiv.quotient_msk\[4\] VSS
+ VSS VCC VCC _0332_ sky130_fd_sc_hs__a22o_1
X_3911_ _1250_ i_op1[9] _1599_ VSS VSS VCC VCC _1607_ sky130_fd_sc_hs__mux2_1
X_3842_ _0672_ _1559_ _1560_ _0800_ VSS VSS VCC VCC _1561_ sky130_fd_sc_hs__o211a_1
X_3773_ _1331_ _1493_ _1495_ _1496_ _0728_ VSS VSS VCC VCC _1497_ sky130_fd_sc_hs__o221a_1
X_5512_ clknet_leaf_50_i_clk _0160_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[30\]
+ sky130_fd_sc_hs__dfxtp_2
X_2724_ u_muldiv.i_op2_signed alu_ctrl\[2\] VSS VSS VCC VCC _0539_ sky130_fd_sc_hs__or2_2
X_2655_ _0469_ VSS VSS VCC VCC _0470_ sky130_fd_sc_hs__clkinv_2
X_5443_ clknet_leaf_2_i_clk _0091_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[3\]
+ sky130_fd_sc_hs__dfxtp_1
X_5374_ clknet_leaf_47_i_clk _0022_ VSS VSS VCC VCC u_bits.i_op1\[6\] sky130_fd_sc_hs__dfxtp_1
X_4325_ _1112_ _1847_ VSS VSS VCC VCC _1848_ sky130_fd_sc_hs__xor2_1
X_4256_ _1802_ VSS VSS VCC VCC _0174_ sky130_fd_sc_hs__clkbuf_1
X_4187_ _1766_ VSS VSS VCC VCC _0141_ sky130_fd_sc_hs__clkbuf_1
X_3207_ _0996_ u_bits.i_op2\[27\] _0636_ _1007_ VSS VSS VCC VCC _1008_ sky130_fd_sc_hs__o22a_1
X_3138_ u_bits.i_op1\[25\] VSS VSS VCC VCC _0943_ sky130_fd_sc_hs__buf_4
X_3069_ _0873_ _0877_ _0524_ VSS VSS VCC VCC _0878_ sky130_fd_sc_hs__mux2_1
Xclkbuf_leaf_52_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_52_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5090_ _2288_ _2437_ VSS VSS VCC VCC _2438_ sky130_fd_sc_hs__nor2_1
X_4110_ u_pc_sel.i_pc_next\[15\] i_pc_next[15] _1723_ VSS VSS VCC VCC _1728_
+ sky130_fd_sc_hs__mux2_1
X_4041_ _1665_ _1684_ _1685_ VSS VSS VCC VCC _0076_ sky130_fd_sc_hs__a21o_1
X_4943_ u_muldiv.on_wait VSS VSS VCC VCC _2303_ sky130_fd_sc_hs__clkbuf_4
X_4874_ u_muldiv.quotient_msk\[29\] _2264_ _2229_ VSS VSS VCC VCC _2269_ sky130_fd_sc_hs__mux2_1
X_3825_ u_bits.i_op2\[17\] _0647_ _0637_ _1544_ VSS VSS VCC VCC _1545_ sky130_fd_sc_hs__o22a_1
X_3756_ u_muldiv.mul\[44\] _0741_ _1480_ VSS VSS VCC VCC _1481_ sky130_fd_sc_hs__a21oi_1
X_2707_ _0500_ _0501_ VSS VSS VCC VCC _0522_ sky130_fd_sc_hs__nand2_1
X_3687_ _1333_ csr_data\[7\] _1388_ VSS VSS VCC VCC _1417_ sky130_fd_sc_hs__o21ai_1
X_5426_ clknet_leaf_52_i_clk _0074_ VSS VSS VCC VCC u_bits.i_op2\[17\] sky130_fd_sc_hs__dfxtp_4
X_2638_ _0452_ VSS VSS VCC VCC _0453_ sky130_fd_sc_hs__clkbuf_4
X_5357_ clknet_leaf_39_i_clk _0005_ VSS VSS VCC VCC u_muldiv.mul\[53\] sky130_fd_sc_hs__dfxtp_1
X_5288_ u_muldiv.divisor\[4\] _2284_ _2285_ u_muldiv.divisor\[5\] VSS VSS VCC
+ VCC _0395_ sky130_fd_sc_hs__a22o_1
X_4308_ _1831_ VSS VSS VCC VCC _1832_ sky130_fd_sc_hs__buf_2
X_4239_ _1793_ VSS VSS VCC VCC _0166_ sky130_fd_sc_hs__clkbuf_1
X_4590_ op_cnt\[0\] op_cnt\[1\] _1204_ VSS VSS VCC VCC _2018_ sky130_fd_sc_hs__a21oi_1
X_3610_ _1343_ _0861_ _0668_ VSS VSS VCC VCC _1344_ sky130_fd_sc_hs__mux2_1
X_3541_ u_muldiv.mul\[0\] _0717_ _0719_ u_muldiv.mul\[32\] _1277_ VSS VSS VCC
+ VCC _1278_ sky130_fd_sc_hs__a221o_1
X_3472_ o_wdata[2] u_wr_mux.i_reg_data2\[18\] _1224_ VSS VSS VCC VCC _1227_
+ sky130_fd_sc_hs__mux2_1
X_5211_ _0904_ _2537_ VSS VSS VCC VCC _2548_ sky130_fd_sc_hs__or2_1
X_5142_ u_muldiv.dividend\[18\] _2484_ _2485_ VSS VSS VCC VCC _2486_ sky130_fd_sc_hs__mux2_1
X_5073_ _2422_ VSS VSS VCC VCC _0371_ sky130_fd_sc_hs__clkbuf_1
X_4024_ _1665_ _1672_ _1673_ VSS VSS VCC VCC _0071_ sky130_fd_sc_hs__a21o_1
X_4926_ u_muldiv.dividend\[0\] u_muldiv.dividend\[1\] VSS VSS VCC VCC _2287_
+ sky130_fd_sc_hs__or2_1
X_4857_ _2161_ _2255_ u_muldiv.o_div\[25\] VSS VSS VCC VCC _2256_ sky130_fd_sc_hs__a21oi_1
X_3808_ _0751_ _1528_ _0712_ VSS VSS VCC VCC _1529_ sky130_fd_sc_hs__o21a_1
X_4788_ u_muldiv.o_div\[11\] _2194_ u_muldiv.o_div\[12\] VSS VSS VCC VCC _2200_
+ sky130_fd_sc_hs__o21ai_1
X_3739_ u_muldiv.dividend\[11\] _1326_ _1327_ u_muldiv.o_div\[11\] _1383_ VSS VSS
+ VCC VCC _1465_ sky130_fd_sc_hs__a221o_1
X_5409_ clknet_leaf_49_i_clk _0057_ VSS VSS VCC VCC u_bits.i_op2\[0\] sky130_fd_sc_hs__dfxtp_1
X_5760_ clknet_leaf_19_i_clk _0403_ VSS VSS VCC VCC u_muldiv.divisor\[12\]
+ sky130_fd_sc_hs__dfxtp_1
X_2972_ u_bits.i_op1\[8\] VSS VSS VCC VCC _0785_ sky130_fd_sc_hs__buf_4
X_5691_ clknet_leaf_26_i_clk _0334_ VSS VSS VCC VCC u_muldiv.quotient_msk\[5\]
+ sky130_fd_sc_hs__dfxtp_1
X_4711_ u_muldiv.divisor\[30\] u_muldiv.dividend\[30\] VSS VSS VCC VCC _2134_
+ sky130_fd_sc_hs__xor2_2
X_4642_ _2060_ u_muldiv.dividend\[2\] _2062_ _2063_ _2064_ VSS VSS VCC VCC
+ _2065_ sky130_fd_sc_hs__a221o_1
X_4573_ o_add[22] _2004_ VSS VSS VCC VCC _2012_ sky130_fd_sc_hs__and2_1
X_3524_ _0653_ _0647_ _0645_ _0646_ _0650_ _0648_ VSS VSS VCC VCC _1261_ sky130_fd_sc_hs__mux4_1
X_3455_ u_wr_mux.i_reg_data2\[10\] o_wdata[2] _0718_ VSS VSS VCC VCC _1218_
+ sky130_fd_sc_hs__mux2_1
X_3386_ _0523_ _0601_ _0608_ _0612_ VSS VSS VCC VCC _1164_ sky130_fd_sc_hs__a31o_1
X_5125_ _0647_ _2293_ _2469_ VSS VSS VCC VCC _2470_ sky130_fd_sc_hs__nand3_1
X_5056_ _2405_ _2406_ _2375_ VSS VSS VCC VCC _2407_ sky130_fd_sc_hs__a21oi_1
X_4007_ _1641_ _1660_ _1661_ VSS VSS VCC VCC _0066_ sky130_fd_sc_hs__a21o_1
X_4909_ u_muldiv.quotient_msk\[18\] _2282_ _2281_ u_muldiv.quotient_msk\[19\] VSS
+ VSS VCC VCC _0347_ sky130_fd_sc_hs__a22o_1
X_3240_ _0747_ _1037_ _1038_ _0453_ VSS VSS VCC VCC _1039_ sky130_fd_sc_hs__a31o_1
X_3171_ _0825_ _0524_ _0840_ VSS VSS VCC VCC _0974_ sky130_fd_sc_hs__and3b_1
X_5743_ clknet_leaf_21_i_clk _0386_ VSS VSS VCC VCC u_muldiv.dividend\[27\]
+ sky130_fd_sc_hs__dfxtp_4
X_2955_ u_bits.i_op1\[21\] VSS VSS VCC VCC _0768_ sky130_fd_sc_hs__buf_4
X_5674_ clknet_leaf_30_i_clk _0317_ VSS VSS VCC VCC u_muldiv.o_div\[20\] sky130_fd_sc_hs__dfxtp_1
X_2886_ _0698_ _0700_ _0663_ VSS VSS VCC VCC _0701_ sky130_fd_sc_hs__mux2_1
X_4625_ u_muldiv.divisor\[10\] u_muldiv.dividend\[10\] VSS VSS VCC VCC _2048_
+ sky130_fd_sc_hs__or2b_1
X_4556_ _1151_ _2006_ VSS VSS VCC VCC _0270_ sky130_fd_sc_hs__nor2_1
X_3507_ _1243_ _1245_ VSS VSS VCC VCC o_wsel[2] sky130_fd_sc_hs__nor2_4
X_4487_ _1974_ VSS VSS VCC VCC _0233_ sky130_fd_sc_hs__clkbuf_1
X_3438_ u_muldiv.i_on_end VSS VSS VCC VCC _1206_ sky130_fd_sc_hs__buf_4
X_3369_ _1151_ VSS VSS VCC VCC o_add[10] sky130_fd_sc_hs__inv_2
X_5108_ _1878_ _2446_ _2454_ VSS VSS VCC VCC _2455_ sky130_fd_sc_hs__o21ai_1
X_5039_ u_muldiv.dividend\[9\] _2391_ _2378_ VSS VSS VCC VCC _2392_ sky130_fd_sc_hs__mux2_1
X_2740_ u_bits.i_op1\[7\] u_muldiv.add_prev\[7\] _0448_ VSS VSS VCC VCC _0555_
+ sky130_fd_sc_hs__mux2_1
X_2671_ _0457_ _0485_ VSS VSS VCC VCC _0486_ sky130_fd_sc_hs__xnor2_1
X_4410_ u_bits.i_op2\[17\] _1915_ VSS VSS VCC VCC _1917_ sky130_fd_sc_hs__or2_1
X_5390_ clknet_leaf_48_i_clk _0038_ VSS VSS VCC VCC u_bits.i_op1\[22\] sky130_fd_sc_hs__dfxtp_2
X_4341_ _0688_ _1859_ _1852_ _1856_ VSS VSS VCC VCC _1861_ sky130_fd_sc_hs__a31o_1
X_4272_ _1810_ VSS VSS VCC VCC _0182_ sky130_fd_sc_hs__clkbuf_1
X_3223_ _1021_ _1022_ VSS VSS VCC VCC _1023_ sky130_fd_sc_hs__and2_1
X_3154_ _0739_ csr_data\[25\] _0958_ _0732_ VSS VSS VCC VCC o_result[25] sky130_fd_sc_hs__o211a_2
X_3085_ _0812_ _0853_ VSS VSS VCC VCC _0893_ sky130_fd_sc_hs__nand2_1
X_3987_ _1641_ _1646_ _1647_ VSS VSS VCC VCC _0060_ sky130_fd_sc_hs__a21o_1
X_5726_ clknet_leaf_20_i_clk _0369_ VSS VSS VCC VCC u_muldiv.dividend\[10\]
+ sky130_fd_sc_hs__dfxtp_2
X_2938_ _0643_ VSS VSS VCC VCC _0751_ sky130_fd_sc_hs__clkbuf_4
X_5657_ clknet_leaf_25_i_clk _0300_ VSS VSS VCC VCC u_muldiv.o_div\[3\] sky130_fd_sc_hs__dfxtp_1
X_2869_ _0672_ _0681_ _0683_ VSS VSS VCC VCC _0684_ sky130_fd_sc_hs__a21oi_1
X_4608_ u_muldiv.divisor\[22\] u_muldiv.dividend\[22\] VSS VSS VCC VCC _2031_
+ sky130_fd_sc_hs__and2b_1
X_5588_ clknet_leaf_23_i_clk _0235_ VSS VSS VCC VCC u_muldiv.mul\[5\] sky130_fd_sc_hs__dfxtp_1
X_4539_ _2001_ VSS VSS VCC VCC _0258_ sky130_fd_sc_hs__clkbuf_1
X_4890_ u_muldiv.quotient_msk\[2\] _1210_ _2279_ u_muldiv.quotient_msk\[3\] VSS
+ VSS VCC VCC _0331_ sky130_fd_sc_hs__a22o_1
X_3910_ _1606_ VSS VSS VCC VCC _0024_ sky130_fd_sc_hs__clkbuf_1
X_3841_ _0687_ _1318_ VSS VSS VCC VCC _1560_ sky130_fd_sc_hs__nand2_1
X_3772_ u_muldiv.mul\[13\] _0748_ _1400_ VSS VSS VCC VCC _1496_ sky130_fd_sc_hs__o21ai_1
X_2723_ _0536_ _0537_ VSS VSS VCC VCC _0538_ sky130_fd_sc_hs__xor2_4
X_5511_ clknet_leaf_49_i_clk _0159_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[29\]
+ sky130_fd_sc_hs__dfxtp_2
X_2654_ _0467_ _0468_ VSS VSS VCC VCC _0469_ sky130_fd_sc_hs__xnor2_1
X_5442_ clknet_leaf_1_i_clk _0090_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[2\]
+ sky130_fd_sc_hs__dfxtp_1
X_5373_ clknet_leaf_47_i_clk _0021_ VSS VSS VCC VCC u_bits.i_op1\[5\] sky130_fd_sc_hs__dfxtp_2
X_4324_ _0831_ _1846_ VSS VSS VCC VCC _1847_ sky130_fd_sc_hs__nand2_1
X_4255_ csr_data\[10\] i_csr_data[10] _1800_ VSS VSS VCC VCC _1802_ sky130_fd_sc_hs__mux2_1
X_4186_ u_wr_mux.i_reg_data2\[11\] i_reg_data2[11] _1756_ VSS VSS VCC VCC
+ _1766_ sky130_fd_sc_hs__mux2_1
X_3206_ _0996_ u_bits.i_op2\[27\] _0867_ VSS VSS VCC VCC _1007_ sky130_fd_sc_hs__a21oi_1
X_3137_ _0644_ _0941_ _0712_ VSS VSS VCC VCC _0942_ sky130_fd_sc_hs__o21a_1
X_3068_ _0875_ _0876_ _0696_ VSS VSS VCC VCC _0877_ sky130_fd_sc_hs__mux2_1
X_5709_ clknet_leaf_31_i_clk _0352_ VSS VSS VCC VCC u_muldiv.quotient_msk\[23\]
+ sky130_fd_sc_hs__dfxtp_1
X_4040_ u_bits.i_op2\[19\] _1663_ _1675_ i_op2[19] VSS VSS VCC VCC _1685_
+ sky130_fd_sc_hs__a22o_1
X_4942_ u_muldiv.dividend\[2\] _2287_ VSS VSS VCC VCC _2302_ sky130_fd_sc_hs__nand2_1
X_4873_ u_muldiv.o_div\[29\] _1835_ _2264_ _2196_ VSS VSS VCC VCC _2268_ sky130_fd_sc_hs__a31o_1
X_3824_ _0618_ _0639_ _1543_ VSS VSS VCC VCC _1544_ sky130_fd_sc_hs__and3_1
X_3755_ u_muldiv.dividend\[12\] _0742_ _0743_ u_muldiv.o_div\[12\] _1383_ VSS VSS
+ VCC VCC _1480_ sky130_fd_sc_hs__a221o_1
X_3686_ _0454_ _1412_ _1414_ _1415_ _1357_ VSS VSS VCC VCC _1416_ sky130_fd_sc_hs__o221a_1
X_2706_ _0515_ _0519_ _0520_ VSS VSS VCC VCC _0521_ sky130_fd_sc_hs__o21a_1
X_5425_ clknet_leaf_52_i_clk _0073_ VSS VSS VCC VCC u_bits.i_op2\[16\] sky130_fd_sc_hs__dfxtp_4
X_2637_ _0451_ VSS VSS VCC VCC _0452_ sky130_fd_sc_hs__buf_4
X_5356_ clknet_leaf_39_i_clk _0004_ VSS VSS VCC VCC u_muldiv.mul\[52\] sky130_fd_sc_hs__dfxtp_1
X_5287_ u_muldiv.divisor\[3\] _2284_ _2285_ u_muldiv.divisor\[4\] VSS VSS VCC
+ VCC _0394_ sky130_fd_sc_hs__a22o_1
X_4307_ _1830_ VSS VSS VCC VCC _1831_ sky130_fd_sc_hs__buf_2
X_4238_ csr_data\[2\] i_csr_data[2] _1789_ VSS VSS VCC VCC _1793_ sky130_fd_sc_hs__mux2_1
X_4169_ _1757_ VSS VSS VCC VCC _0132_ sky130_fd_sc_hs__clkbuf_1
X_3540_ u_muldiv.dividend\[0\] _0633_ _0722_ u_muldiv.o_div\[0\] VSS VSS VCC
+ VCC _1277_ sky130_fd_sc_hs__a22o_1
X_5210_ _2109_ _2546_ VSS VSS VCC VCC _2547_ sky130_fd_sc_hs__xnor2_1
X_3471_ _1226_ VSS VSS VCC VCC o_wdata[17] sky130_fd_sc_hs__buf_2
X_5141_ _2153_ VSS VSS VCC VCC _2485_ sky130_fd_sc_hs__buf_4
X_5072_ u_muldiv.dividend\[12\] _2421_ _2378_ VSS VSS VCC VCC _2422_ sky130_fd_sc_hs__mux2_1
X_4023_ u_bits.i_op2\[14\] _1663_ _1651_ i_op2[14] VSS VSS VCC VCC _1673_
+ sky130_fd_sc_hs__a22o_1
X_4925_ u_muldiv.dividend\[0\] u_muldiv.dividend\[1\] VSS VSS VCC VCC _2286_
+ sky130_fd_sc_hs__nand2_1
X_4856_ u_muldiv.quotient_msk\[25\] _2250_ _2229_ VSS VSS VCC VCC _2255_ sky130_fd_sc_hs__mux2_1
X_3807_ _0910_ _1262_ _0879_ VSS VSS VCC VCC _1528_ sky130_fd_sc_hs__mux2_1
X_4787_ _2181_ _2197_ _2199_ VSS VSS VCC VCC _0308_ sky130_fd_sc_hs__a21oi_1
Xclkbuf_leaf_51_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_51_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3738_ _0714_ _1462_ _1463_ _0623_ _1150_ VSS VSS VCC VCC _1464_ sky130_fd_sc_hs__o32a_1
X_3669_ _0453_ VSS VSS VCC VCC _1400_ sky130_fd_sc_hs__clkbuf_2
X_5408_ clknet_leaf_1_i_clk _0056_ VSS VSS VCC VCC u_pc_sel.i_inst_branch
+ sky130_fd_sc_hs__dfxtp_1
X_5339_ _1141_ _1585_ VSS VSS VCC VCC _0432_ sky130_fd_sc_hs__nor2_1
Xclkbuf_leaf_19_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_19_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_2971_ _0781_ _0782_ _0783_ VSS VSS VCC VCC _0784_ sky130_fd_sc_hs__mux2_2
X_5690_ clknet_leaf_26_i_clk _0333_ VSS VSS VCC VCC u_muldiv.quotient_msk\[4\]
+ sky130_fd_sc_hs__dfxtp_1
X_4710_ u_muldiv.dividend\[29\] u_muldiv.divisor\[29\] VSS VSS VCC VCC _2133_
+ sky130_fd_sc_hs__and2b_1
X_4641_ u_muldiv.divisor\[1\] u_muldiv.dividend\[1\] VSS VSS VCC VCC _2064_
+ sky130_fd_sc_hs__and2b_1
X_4572_ _2011_ VSS VSS VCC VCC _0281_ sky130_fd_sc_hs__clkbuf_1
X_3523_ _1256_ _1259_ _0789_ VSS VSS VCC VCC _1260_ sky130_fd_sc_hs__mux2_1
X_3454_ _1217_ VSS VSS VCC VCC o_wdata[9] sky130_fd_sc_hs__buf_2
X_3385_ _1163_ VSS VSS VCC VCC o_add[14] sky130_fd_sc_hs__inv_2
X_5124_ u_bits.i_op1\[15\] u_bits.i_op1\[16\] _2450_ VSS VSS VCC VCC _2469_
+ sky130_fd_sc_hs__or3_2
X_5055_ _2047_ _2078_ VSS VSS VCC VCC _2406_ sky130_fd_sc_hs__and2b_1
X_4006_ u_bits.i_op2\[9\] _1637_ _1651_ i_op2[9] VSS VSS VCC VCC _1661_ sky130_fd_sc_hs__a22o_1
X_4908_ u_muldiv.quotient_msk\[17\] _2282_ _2281_ u_muldiv.quotient_msk\[18\] VSS
+ VSS VCC VCC _0346_ sky130_fd_sc_hs__a22o_1
X_4839_ u_muldiv.o_div\[21\] u_muldiv.o_div\[22\] _2233_ VSS VSS VCC VCC _2241_
+ sky130_fd_sc_hs__or3_2
X_3170_ _0836_ _0838_ _0760_ VSS VSS VCC VCC _0973_ sky130_fd_sc_hs__mux2_1
X_5742_ clknet_leaf_21_i_clk _0385_ VSS VSS VCC VCC u_muldiv.dividend\[26\]
+ sky130_fd_sc_hs__dfxtp_4
X_2954_ _0751_ _0766_ _0712_ VSS VSS VCC VCC _0767_ sky130_fd_sc_hs__o21a_1
X_5673_ clknet_leaf_30_i_clk _0316_ VSS VSS VCC VCC u_muldiv.o_div\[19\] sky130_fd_sc_hs__dfxtp_1
X_2885_ _0699_ u_bits.i_op1\[31\] _0649_ VSS VSS VCC VCC _0700_ sky130_fd_sc_hs__mux2_1
X_4624_ u_muldiv.dividend\[11\] u_muldiv.divisor\[11\] VSS VSS VCC VCC _2047_
+ sky130_fd_sc_hs__and2b_1
X_4555_ _1145_ _2006_ VSS VSS VCC VCC _0269_ sky130_fd_sc_hs__nor2_1
X_3506_ _1224_ o_add[1] VSS VSS VCC VCC _1245_ sky130_fd_sc_hs__nor2_2
X_4486_ u_muldiv.mul\[3\] u_muldiv.mul\[4\] _1584_ VSS VSS VCC VCC _1974_
+ sky130_fd_sc_hs__mux2_1
X_3437_ i_alu_ctrl[1] VSS VSS VCC VCC _1205_ sky130_fd_sc_hs__inv_2
X_3368_ _0589_ _1148_ VSS VSS VCC VCC _1151_ sky130_fd_sc_hs__xnor2_4
X_5107_ _2303_ _2449_ _2453_ _1829_ VSS VSS VCC VCC _2454_ sky130_fd_sc_hs__a22o_1
X_3299_ _0739_ csr_data\[30\] _1093_ _0732_ VSS VSS VCC VCC o_result[30] sky130_fd_sc_hs__o211a_2
X_5038_ _1208_ _2380_ _2381_ _2390_ VSS VSS VCC VCC _2391_ sky130_fd_sc_hs__a31o_1
X_2670_ _0460_ u_bits.i_op2\[17\] u_bits.i_op1\[17\] _0464_ VSS VSS VCC VCC
+ _0485_ sky130_fd_sc_hs__a22o_1
X_4340_ _1859_ _1850_ _0688_ VSS VSS VCC VCC _1860_ sky130_fd_sc_hs__a21oi_1
X_4271_ csr_data\[18\] i_csr_data[18] _1800_ VSS VSS VCC VCC _1810_ sky130_fd_sc_hs__mux2_1
X_3222_ _1019_ _1020_ VSS VSS VCC VCC _1022_ sky130_fd_sc_hs__or2_1
X_3153_ _0939_ _0957_ _0447_ VSS VSS VCC VCC _0958_ sky130_fd_sc_hs__a21o_1
X_3084_ u_muldiv.mul\[24\] _0740_ _0741_ u_muldiv.mul\[56\] _0891_ VSS VSS VCC
+ VCC _0892_ sky130_fd_sc_hs__a221o_1
X_3986_ _0909_ _1637_ _1638_ i_op2[3] VSS VSS VCC VCC _1647_ sky130_fd_sc_hs__a22o_1
X_5725_ clknet_leaf_26_i_clk _0368_ VSS VSS VCC VCC u_muldiv.dividend\[9\]
+ sky130_fd_sc_hs__dfxtp_1
X_2937_ _0749_ VSS VSS VCC VCC _0750_ sky130_fd_sc_hs__buf_2
X_5656_ clknet_leaf_24_i_clk _0299_ VSS VSS VCC VCC u_muldiv.o_div\[2\] sky130_fd_sc_hs__dfxtp_1
X_4607_ u_muldiv.divisor\[28\] u_muldiv.dividend\[28\] VSS VSS VCC VCC _2030_
+ sky130_fd_sc_hs__nand2b_4
X_2868_ _0625_ _0682_ VSS VSS VCC VCC _0683_ sky130_fd_sc_hs__nand2_1
X_5587_ clknet_leaf_23_i_clk _0234_ VSS VSS VCC VCC u_muldiv.mul\[4\] sky130_fd_sc_hs__dfxtp_1
X_2799_ _0523_ _0601_ _0608_ _0613_ _0484_ VSS VSS VCC VCC _0614_ sky130_fd_sc_hs__a311o_1
X_4538_ u_muldiv.mul\[28\] u_muldiv.mul\[29\] _1583_ VSS VSS VCC VCC _2001_
+ sky130_fd_sc_hs__mux2_1
X_4469_ u_bits.i_op2\[29\] _1852_ _1962_ _1831_ VSS VSS VCC VCC _1964_ sky130_fd_sc_hs__a31o_1
X_3840_ _0833_ _0835_ _0836_ _0838_ _0825_ _0707_ VSS VSS VCC VCC _1559_ sky130_fd_sc_hs__mux4_1
X_3771_ u_muldiv.mul\[45\] _0741_ _1494_ VSS VSS VCC VCC _1495_ sky130_fd_sc_hs__a21oi_1
X_2722_ u_bits.i_op1\[1\] u_muldiv.add_prev\[1\] _0449_ VSS VSS VCC VCC _0537_
+ sky130_fd_sc_hs__mux2_2
X_5510_ clknet_leaf_49_i_clk _0158_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[28\]
+ sky130_fd_sc_hs__dfxtp_2
X_2653_ u_bits.i_op1\[20\] u_muldiv.add_prev\[20\] _0451_ VSS VSS VCC VCC
+ _0468_ sky130_fd_sc_hs__mux2_1
X_5441_ clknet_leaf_1_i_clk _0089_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[1\]
+ sky130_fd_sc_hs__dfxtp_1
X_5372_ clknet_leaf_47_i_clk _0020_ VSS VSS VCC VCC u_bits.i_op1\[4\] sky130_fd_sc_hs__dfxtp_2
X_4323_ _1845_ VSS VSS VCC VCC _1846_ sky130_fd_sc_hs__buf_2
X_4254_ _1801_ VSS VSS VCC VCC _0173_ sky130_fd_sc_hs__clkbuf_1
X_4185_ _1765_ VSS VSS VCC VCC _0140_ sky130_fd_sc_hs__clkbuf_1
X_3205_ _0674_ _1004_ _1005_ VSS VSS VCC VCC _1006_ sky130_fd_sc_hs__a21o_1
X_3136_ _0909_ _0940_ _0911_ VSS VSS VCC VCC _0941_ sky130_fd_sc_hs__o21a_1
X_3067_ u_bits.i_op1\[11\] u_bits.i_op1\[10\] u_bits.i_op1\[9\] u_bits.i_op1\[8\]
+ _0657_ _0663_ VSS VSS VCC VCC _0876_ sky130_fd_sc_hs__mux4_1
X_5708_ clknet_leaf_30_i_clk _0351_ VSS VSS VCC VCC u_muldiv.quotient_msk\[22\]
+ sky130_fd_sc_hs__dfxtp_1
X_3969_ i_rd[3] _1632_ _1636_ o_rd[3] VSS VSS VCC VCC _0053_ sky130_fd_sc_hs__a22o_1
X_5639_ clknet_leaf_41_i_clk _0286_ VSS VSS VCC VCC u_muldiv.add_prev\[25\]
+ sky130_fd_sc_hs__dfxtp_1
X_4941_ u_muldiv.dividend\[0\] u_muldiv.dividend\[1\] u_muldiv.dividend\[2\] VSS
+ VSS VCC VCC _2301_ sky130_fd_sc_hs__or3_1
X_4872_ _2267_ VSS VSS VCC VCC _0325_ sky130_fd_sc_hs__clkbuf_1
X_3823_ u_bits.i_op2\[17\] _0647_ VSS VSS VCC VCC _1543_ sky130_fd_sc_hs__nand2_1
X_3754_ _0714_ _1477_ _1478_ _0623_ _1157_ VSS VSS VCC VCC _1479_ sky130_fd_sc_hs__o32a_1
X_3685_ u_muldiv.mul\[7\] _1330_ _1400_ VSS VSS VCC VCC _1415_ sky130_fd_sc_hs__o21ai_1
X_2705_ _0513_ _0514_ VSS VSS VCC VCC _0520_ sky130_fd_sc_hs__nand2_1
X_2636_ _0450_ VSS VSS VCC VCC _0451_ sky130_fd_sc_hs__clkbuf_4
X_5424_ clknet_leaf_52_i_clk _0072_ VSS VSS VCC VCC u_bits.i_op2\[15\] sky130_fd_sc_hs__dfxtp_4
X_5355_ _0616_ _2004_ VSS VSS VCC VCC _0445_ sky130_fd_sc_hs__nor2_1
X_5286_ u_muldiv.divisor\[2\] _2284_ _2285_ u_muldiv.divisor\[3\] VSS VSS VCC
+ VCC _0393_ sky130_fd_sc_hs__a22o_1
X_4306_ u_muldiv.on_wait u_muldiv.i_on_end VSS VSS VCC VCC _1830_ sky130_fd_sc_hs__or2_1
X_4237_ _1792_ VSS VSS VCC VCC _0165_ sky130_fd_sc_hs__clkbuf_1
X_4168_ o_wdata[2] i_reg_data2[2] _1756_ VSS VSS VCC VCC _1757_ sky130_fd_sc_hs__mux2_1
X_4099_ u_pc_sel.i_pc_next\[10\] i_pc_next[10] _1712_ VSS VSS VCC VCC _1722_
+ sky130_fd_sc_hs__mux2_1
X_3119_ _0636_ VSS VSS VCC VCC _0926_ sky130_fd_sc_hs__clkbuf_4
X_3470_ o_wdata[1] u_wr_mux.i_reg_data2\[17\] _1224_ VSS VSS VCC VCC _1226_
+ sky130_fd_sc_hs__mux2_1
X_5140_ _2476_ _2483_ _1877_ VSS VSS VCC VCC _2484_ sky130_fd_sc_hs__mux2_1
X_5071_ _2414_ _2420_ _1877_ VSS VSS VCC VCC _2421_ sky130_fd_sc_hs__mux2_1
X_4022_ u_bits.i_op2\[15\] _1487_ _1657_ VSS VSS VCC VCC _1672_ sky130_fd_sc_hs__mux2_1
X_4924_ u_muldiv.quotient_msk\[30\] _2284_ _2285_ u_muldiv.quotient_msk\[31\] VSS
+ VSS VCC VCC _0359_ sky130_fd_sc_hs__a22o_1
X_4855_ u_muldiv.o_div\[25\] _2170_ _2250_ _2196_ VSS VSS VCC VCC _2254_ sky130_fd_sc_hs__a31o_1
X_4786_ _2167_ _2198_ u_muldiv.o_div\[11\] VSS VSS VCC VCC _2199_ sky130_fd_sc_hs__a21oi_1
X_3806_ u_muldiv.mul\[16\] _0717_ _0720_ u_muldiv.mul\[48\] _1526_ VSS VSS VCC
+ VCC _1527_ sky130_fd_sc_hs__a221o_1
X_3737_ u_bits.i_op2\[11\] _1251_ _0906_ VSS VSS VCC VCC _1463_ sky130_fd_sc_hs__a21oi_1
X_3668_ u_muldiv.mul\[38\] _1325_ _1398_ VSS VSS VCC VCC _1399_ sky130_fd_sc_hs__a21oi_1
X_3599_ _0454_ _1324_ _1329_ _1332_ _1333_ VSS VSS VCC VCC _1334_ sky130_fd_sc_hs__o221a_1
X_5407_ clknet_leaf_1_i_clk _0055_ VSS VSS VCC VCC u_pc_sel.i_inst_jal_jalr
+ sky130_fd_sc_hs__dfxtp_1
X_5338_ _1142_ _1585_ VSS VSS VCC VCC _0431_ sky130_fd_sc_hs__nor2_1
X_5269_ u_muldiv.dividend\[30\] _2583_ VSS VSS VCC VCC _2601_ sky130_fd_sc_hs__nor2_1
X_2970_ _0663_ VSS VSS VCC VCC _0783_ sky130_fd_sc_hs__clkbuf_4
X_4640_ u_muldiv.dividend\[0\] u_muldiv.divisor\[0\] VSS VSS VCC VCC _2063_
+ sky130_fd_sc_hs__or2b_1
X_4571_ o_add[21] _2004_ VSS VSS VCC VCC _2011_ sky130_fd_sc_hs__and2_1
X_3522_ u_bits.i_op1\[4\] _1257_ _0786_ _1258_ _0651_ _0783_ VSS VSS VCC VCC
+ _1259_ sky130_fd_sc_hs__mux4_1
X_3453_ u_wr_mux.i_reg_data2\[9\] o_wdata[1] _0718_ VSS VSS VCC VCC _1217_
+ sky130_fd_sc_hs__mux2_1
X_5123_ u_muldiv.dividend\[17\] u_muldiv.dividend\[16\] _2444_ VSS VSS VCC VCC
+ _2468_ sky130_fd_sc_hs__or3_2
X_3384_ _0509_ _1160_ VSS VSS VCC VCC _1163_ sky130_fd_sc_hs__xor2_4
X_5054_ _2048_ _2397_ VSS VSS VCC VCC _2405_ sky130_fd_sc_hs__and2_1
X_4005_ _1445_ u_bits.i_op2\[8\] _1657_ VSS VSS VCC VCC _1660_ sky130_fd_sc_hs__mux2_1
X_4907_ _1209_ VSS VSS VCC VCC _2282_ sky130_fd_sc_hs__buf_2
X_4838_ u_muldiv.o_div\[21\] _2233_ u_muldiv.o_div\[22\] VSS VSS VCC VCC _2240_
+ sky130_fd_sc_hs__o21ai_1
X_4769_ u_muldiv.o_div\[7\] _2179_ u_muldiv.o_div\[8\] VSS VSS VCC VCC _2185_
+ sky130_fd_sc_hs__o21ai_1
Xclkbuf_leaf_50_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_50_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5741_ clknet_leaf_21_i_clk _0384_ VSS VSS VCC VCC u_muldiv.dividend\[25\]
+ sky130_fd_sc_hs__dfxtp_2
X_2953_ _0759_ _0765_ _0707_ VSS VSS VCC VCC _0766_ sky130_fd_sc_hs__mux2_1
X_5672_ clknet_leaf_28_i_clk _0315_ VSS VSS VCC VCC u_muldiv.o_div\[18\] sky130_fd_sc_hs__dfxtp_1
X_2884_ u_bits.i_op1\[30\] VSS VSS VCC VCC _0699_ sky130_fd_sc_hs__clkbuf_4
X_4623_ _2044_ _2045_ VSS VSS VCC VCC _2046_ sky130_fd_sc_hs__nand2_1
X_4554_ _1147_ _2006_ VSS VSS VCC VCC _0268_ sky130_fd_sc_hs__nor2_1
X_3505_ _1242_ _1244_ VSS VSS VCC VCC o_wsel[1] sky130_fd_sc_hs__nor2_4
X_4485_ _1973_ VSS VSS VCC VCC _0232_ sky130_fd_sc_hs__clkbuf_1
X_3436_ _1204_ _1192_ _1203_ VSS VSS VCC VCC mul_op2_signed_next sky130_fd_sc_hs__nor3_1
X_3367_ _1150_ VSS VSS VCC VCC o_add[11] sky130_fd_sc_hs__inv_2
X_5106_ _1206_ _2451_ _2452_ VSS VSS VCC VCC _2453_ sky130_fd_sc_hs__or3_1
X_5037_ _2303_ _2384_ _2389_ VSS VSS VCC VCC _2390_ sky130_fd_sc_hs__a21oi_1
X_3298_ _1079_ _1092_ _0446_ VSS VSS VCC VCC _1093_ sky130_fd_sc_hs__a21o_1
Xclkbuf_leaf_18_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_18_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4270_ _1809_ VSS VSS VCC VCC _0181_ sky130_fd_sc_hs__clkbuf_1
X_3221_ _1019_ _1020_ VSS VSS VCC VCC _1021_ sky130_fd_sc_hs__nand2_1
X_3152_ _0750_ o_add[25] _0954_ _0956_ _0804_ VSS VSS VCC VCC _0957_ sky130_fd_sc_hs__a221o_1
X_3083_ u_muldiv.dividend\[24\] _0742_ _0743_ u_muldiv.o_div\[24\] _0744_ VSS VSS
+ VCC VCC _0891_ sky130_fd_sc_hs__a221o_1
X_3985_ _0688_ _0923_ _1639_ VSS VSS VCC VCC _1646_ sky130_fd_sc_hs__mux2_1
X_5724_ clknet_leaf_26_i_clk _0367_ VSS VSS VCC VCC u_muldiv.dividend\[8\]
+ sky130_fd_sc_hs__dfxtp_2
X_2936_ _0747_ _0748_ VSS VSS VCC VCC _0749_ sky130_fd_sc_hs__nand2_2
X_5655_ clknet_leaf_31_i_clk _0298_ VSS VSS VCC VCC u_muldiv.o_div\[1\] sky130_fd_sc_hs__dfxtp_1
X_2867_ o_funct3[1] o_funct3[0] VSS VSS VCC VCC _0682_ sky130_fd_sc_hs__and2b_1
X_4606_ _1835_ _2026_ _2027_ _2028_ VSS VSS VCC VCC _2029_ sky130_fd_sc_hs__a31o_1
X_5586_ clknet_leaf_23_i_clk _0233_ VSS VSS VCC VCC u_muldiv.mul\[3\] sky130_fd_sc_hs__dfxtp_1
X_2798_ _0610_ _0612_ VSS VSS VCC VCC _0613_ sky130_fd_sc_hs__or2_1
X_4537_ _2000_ VSS VSS VCC VCC _0257_ sky130_fd_sc_hs__clkbuf_1
X_4468_ _1850_ _1962_ u_bits.i_op2\[29\] VSS VSS VCC VCC _1963_ sky130_fd_sc_hs__a21oi_1
X_3419_ _1171_ _1188_ _0618_ VSS VSS VCC VCC _1190_ sky130_fd_sc_hs__a21oi_1
X_4399_ u_bits.i_op2\[15\] _1852_ _1906_ _1856_ VSS VSS VCC VCC _1908_ sky130_fd_sc_hs__a31o_1
X_3770_ u_muldiv.dividend\[13\] _0742_ _0743_ u_muldiv.o_div\[13\] _1383_ VSS VSS
+ VCC VCC _1494_ sky130_fd_sc_hs__a221o_1
X_2721_ _0456_ _0535_ VSS VSS VCC VCC _0536_ sky130_fd_sc_hs__xnor2_2
X_5440_ clknet_leaf_0_i_clk _0088_ VSS VSS VCC VCC u_bits.i_op2\[31\] sky130_fd_sc_hs__dfxtp_4
X_2652_ _0458_ _0466_ VSS VSS VCC VCC _0467_ sky130_fd_sc_hs__xnor2_2
X_5371_ clknet_leaf_46_i_clk _0019_ VSS VSS VCC VCC u_bits.i_op1\[3\] sky130_fd_sc_hs__dfxtp_2
X_4322_ _1844_ VSS VSS VCC VCC _1845_ sky130_fd_sc_hs__buf_2
X_4253_ csr_data\[9\] i_csr_data[9] _1800_ VSS VSS VCC VCC _1801_ sky130_fd_sc_hs__mux2_1
X_3204_ _0669_ _0788_ _0881_ VSS VSS VCC VCC _1005_ sky130_fd_sc_hs__and3b_1
X_4184_ u_wr_mux.i_reg_data2\[10\] i_reg_data2[10] _1756_ VSS VSS VCC VCC
+ _1765_ sky130_fd_sc_hs__mux2_1
X_3135_ _0757_ _0764_ _0696_ VSS VSS VCC VCC _0940_ sky130_fd_sc_hs__mux2_1
X_3066_ _0782_ _0874_ _0533_ VSS VSS VCC VCC _0875_ sky130_fd_sc_hs__mux2_1
X_3968_ i_rd[2] _1632_ _1636_ o_rd[2] VSS VSS VCC VCC _0052_ sky130_fd_sc_hs__a22o_1
X_5707_ clknet_leaf_30_i_clk _0350_ VSS VSS VCC VCC u_muldiv.quotient_msk\[21\]
+ sky130_fd_sc_hs__dfxtp_1
X_2919_ _0461_ u_bits.i_op2\[21\] _0465_ u_bits.i_op1\[21\] VSS VSS VCC VCC
+ _0733_ sky130_fd_sc_hs__a22o_1
X_3899_ _0794_ i_op1[3] _1599_ VSS VSS VCC VCC _1601_ sky130_fd_sc_hs__mux2_1
X_5638_ clknet_leaf_41_i_clk _0285_ VSS VSS VCC VCC u_muldiv.add_prev\[24\]
+ sky130_fd_sc_hs__dfxtp_1
X_5569_ clknet_leaf_9_i_clk _0216_ VSS VSS VCC VCC u_muldiv.divisor\[50\]
+ sky130_fd_sc_hs__dfxtp_1
X_4940_ _2300_ VSS VSS VCC VCC _0360_ sky130_fd_sc_hs__clkbuf_1
X_4871_ u_muldiv.o_div\[28\] _2266_ _2244_ VSS VSS VCC VCC _2267_ sky130_fd_sc_hs__mux2_1
X_3822_ _0751_ _1290_ _0711_ VSS VSS VCC VCC _1542_ sky130_fd_sc_hs__o21a_1
X_3753_ u_bits.i_op2\[12\] _0777_ _0906_ VSS VSS VCC VCC _1478_ sky130_fd_sc_hs__a21oi_1
X_3684_ u_muldiv.mul\[39\] _1325_ _1413_ VSS VSS VCC VCC _1414_ sky130_fd_sc_hs__a21oi_1
X_2704_ _0517_ _0518_ VSS VSS VCC VCC _0519_ sky130_fd_sc_hs__nand2_1
X_2635_ _0449_ VSS VSS VCC VCC _0450_ sky130_fd_sc_hs__buf_4
X_5423_ clknet_leaf_52_i_clk _0071_ VSS VSS VCC VCC u_bits.i_op2\[14\] sky130_fd_sc_hs__dfxtp_4
X_5354_ _2630_ VSS VSS VCC VCC _0444_ sky130_fd_sc_hs__clkbuf_1
X_4305_ _1828_ VSS VSS VCC VCC _1829_ sky130_fd_sc_hs__clkbuf_4
X_5285_ u_muldiv.divisor\[1\] _2284_ _2285_ u_muldiv.divisor\[2\] VSS VSS VCC
+ VCC _0392_ sky130_fd_sc_hs__a22o_1
X_4236_ csr_data\[1\] i_csr_data[1] _1789_ VSS VSS VCC VCC _1792_ sky130_fd_sc_hs__mux2_1
X_4167_ _1711_ VSS VSS VCC VCC _1756_ sky130_fd_sc_hs__clkbuf_4
X_3118_ _0642_ _0683_ VSS VSS VCC VCC _0925_ sky130_fd_sc_hs__nor2_4
X_4098_ _1721_ VSS VSS VCC VCC _0097_ sky130_fd_sc_hs__clkbuf_1
X_3049_ _0627_ VSS VSS VCC VCC _0858_ sky130_fd_sc_hs__buf_2
X_5070_ _1826_ _2415_ _2416_ _2418_ _2419_ VSS VSS VCC VCC _2420_ sky130_fd_sc_hs__a32o_1
X_4021_ _1665_ _1670_ _1671_ VSS VSS VCC VCC _0070_ sky130_fd_sc_hs__a21o_1
X_4923_ _1946_ VSS VSS VCC VCC _2285_ sky130_fd_sc_hs__clkbuf_4
X_4854_ _2253_ VSS VSS VCC VCC _0321_ sky130_fd_sc_hs__clkbuf_1
X_4785_ u_muldiv.quotient_msk\[11\] _2194_ _2156_ VSS VSS VCC VCC _2198_ sky130_fd_sc_hs__mux2_1
X_3805_ u_muldiv.dividend\[16\] _0721_ _0723_ u_muldiv.o_div\[16\] _0724_ VSS VSS
+ VCC VCC _1526_ sky130_fd_sc_hs__a221o_1
X_3736_ _0908_ _1461_ VSS VSS VCC VCC _1462_ sky130_fd_sc_hs__nor2_1
X_3667_ u_muldiv.dividend\[6\] _1326_ _1327_ u_muldiv.o_div\[6\] _1383_ VSS VSS
+ VCC VCC _1398_ sky130_fd_sc_hs__a221o_1
X_3598_ _0728_ VSS VSS VCC VCC _1333_ sky130_fd_sc_hs__buf_2
X_5406_ clknet_leaf_51_i_clk _0054_ VSS VSS VCC VCC o_rd[4] sky130_fd_sc_hs__dfxtp_2
X_5337_ _1135_ _1585_ VSS VSS VCC VCC _0430_ sky130_fd_sc_hs__nor2_1
X_5268_ _2375_ _2595_ _2596_ _2597_ _2599_ VSS VSS VCC VCC _2600_ sky130_fd_sc_hs__a32o_1
X_4219_ _1783_ VSS VSS VCC VCC _0156_ sky130_fd_sc_hs__clkbuf_1
X_5199_ u_bits.i_op1\[21\] _0691_ _0692_ _2511_ VSS VSS VCC VCC _2537_ sky130_fd_sc_hs__or4_2
X_4570_ _0616_ _2007_ VSS VSS VCC VCC _0280_ sky130_fd_sc_hs__nor2_1
X_3521_ u_bits.i_op1\[7\] VSS VSS VCC VCC _1258_ sky130_fd_sc_hs__clkbuf_4
X_3452_ _1216_ VSS VSS VCC VCC o_wdata[8] sky130_fd_sc_hs__buf_2
X_3383_ _1162_ VSS VSS VCC VCC o_add[15] sky130_fd_sc_hs__inv_2
X_5122_ u_muldiv.dividend\[16\] _2444_ u_muldiv.dividend\[17\] VSS VSS VCC VCC
+ _2467_ sky130_fd_sc_hs__o21ai_1
X_5053_ u_muldiv.dividend\[10\] _2380_ u_muldiv.dividend\[11\] VSS VSS VCC VCC
+ _2404_ sky130_fd_sc_hs__o21ai_1
X_4004_ _1641_ _1658_ _1659_ VSS VSS VCC VCC _0065_ sky130_fd_sc_hs__a21o_1
X_4906_ u_muldiv.quotient_msk\[16\] _2280_ _2281_ u_muldiv.quotient_msk\[17\] VSS
+ VSS VCC VCC _0345_ sky130_fd_sc_hs__a22o_1
X_4837_ _2181_ _2237_ _2239_ VSS VSS VCC VCC _0318_ sky130_fd_sc_hs__a21oi_1
X_4768_ _2181_ _2182_ _2184_ VSS VSS VCC VCC _0304_ sky130_fd_sc_hs__a21oi_1
X_4699_ _2031_ _2105_ _2106_ _2119_ _2121_ VSS VSS VCC VCC _2122_ sky130_fd_sc_hs__o311a_1
X_3719_ _1445_ _1305_ _1267_ VSS VSS VCC VCC _1446_ sky130_fd_sc_hs__a21oi_1
X_5740_ clknet_leaf_17_i_clk _0383_ VSS VSS VCC VCC u_muldiv.dividend\[24\]
+ sky130_fd_sc_hs__dfxtp_4
X_2952_ _0760_ _0764_ _0704_ VSS VSS VCC VCC _0765_ sky130_fd_sc_hs__o21a_1
X_5671_ clknet_leaf_31_i_clk _0314_ VSS VSS VCC VCC u_muldiv.o_div\[17\] sky130_fd_sc_hs__dfxtp_1
X_2883_ u_bits.i_op1\[28\] _0697_ _0649_ VSS VSS VCC VCC _0698_ sky130_fd_sc_hs__mux2_1
X_4622_ u_muldiv.dividend\[12\] u_muldiv.divisor\[12\] VSS VSS VCC VCC _2045_
+ sky130_fd_sc_hs__or2b_1
X_4553_ _1141_ _2006_ VSS VSS VCC VCC _0267_ sky130_fd_sc_hs__nor2_1
X_4484_ u_muldiv.mul\[2\] u_muldiv.mul\[3\] _1584_ VSS VSS VCC VCC _1973_
+ sky130_fd_sc_hs__mux2_1
X_3504_ _0621_ o_add[0] VSS VSS VCC VCC _1244_ sky130_fd_sc_hs__nor2_2
X_3435_ o_ready VSS VSS VCC VCC _1204_ sky130_fd_sc_hs__clkbuf_4
X_3366_ _0584_ _1149_ VSS VSS VCC VCC _1150_ sky130_fd_sc_hs__xnor2_4
X_5105_ _2293_ _2450_ _0654_ VSS VSS VCC VCC _2452_ sky130_fd_sc_hs__a21oi_1
X_3297_ _0750_ o_add[30] _1090_ _1091_ _0804_ VSS VSS VCC VCC _1092_ sky130_fd_sc_hs__a221o_1
X_5036_ _1206_ _2387_ _2388_ _1828_ VSS VSS VCC VCC _2389_ sky130_fd_sc_hs__o31a_1
X_3220_ u_bits.i_op1\[28\] u_muldiv.add_prev\[28\] _0452_ VSS VSS VCC VCC
+ _1020_ sky130_fd_sc_hs__mux2_1
X_3151_ _0629_ _0950_ _0955_ VSS VSS VCC VCC _0956_ sky130_fd_sc_hs__a21oi_1
X_3082_ _0739_ csr_data\[23\] _0890_ VSS VSS VCC VCC o_result[23] sky130_fd_sc_hs__o21a_2
X_3984_ _1641_ _1644_ _1645_ VSS VSS VCC VCC _0059_ sky130_fd_sc_hs__a21o_1
X_5723_ clknet_leaf_26_i_clk _0366_ VSS VSS VCC VCC u_muldiv.dividend\[7\]
+ sky130_fd_sc_hs__dfxtp_1
X_2935_ _0625_ _0639_ VSS VSS VCC VCC _0748_ sky130_fd_sc_hs__nand2_2
X_5654_ clknet_leaf_22_i_clk u_muldiv.i_on_wait VSS VSS VCC VCC u_muldiv.on_wait
+ sky130_fd_sc_hs__dfxtp_2
X_2866_ _0674_ _0680_ VSS VSS VCC VCC _0681_ sky130_fd_sc_hs__nand2_1
X_4605_ u_muldiv.quotient_msk\[1\] u_muldiv.o_div\[1\] _1841_ VSS VSS VCC VCC
+ _2028_ sky130_fd_sc_hs__o21a_1
X_5585_ clknet_leaf_23_i_clk _0232_ VSS VSS VCC VCC u_muldiv.mul\[2\] sky130_fd_sc_hs__dfxtp_1
X_2797_ _0492_ _0611_ VSS VSS VCC VCC _0612_ sky130_fd_sc_hs__nand2_2
X_4536_ u_muldiv.mul\[27\] u_muldiv.mul\[28\] _1989_ VSS VSS VCC VCC _2000_
+ sky130_fd_sc_hs__mux2_1
X_4467_ u_bits.i_op2\[28\] _1958_ VSS VSS VCC VCC _1962_ sky130_fd_sc_hs__or2_1
X_4398_ _1868_ _1906_ u_bits.i_op2\[15\] VSS VSS VCC VCC _1907_ sky130_fd_sc_hs__a21oi_1
X_3418_ _1171_ _1188_ VSS VSS VCC VCC _1189_ sky130_fd_sc_hs__or2_1
X_3349_ _1137_ VSS VSS VCC VCC o_add[4] sky130_fd_sc_hs__inv_2
X_5019_ _1258_ _2363_ _2293_ VSS VSS VCC VCC _2373_ sky130_fd_sc_hs__o21ai_1
X_2720_ _0448_ u_bits.i_op1\[1\] _0497_ _0534_ VSS VSS VCC VCC _0535_ sky130_fd_sc_hs__a31o_1
X_2651_ _0461_ u_bits.i_op2\[20\] _0465_ u_bits.i_op1\[20\] VSS VSS VCC VCC
+ _0466_ sky130_fd_sc_hs__a22o_1
Xclkbuf_leaf_17_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_17_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5370_ clknet_leaf_47_i_clk _0018_ VSS VSS VCC VCC u_bits.i_op1\[2\] sky130_fd_sc_hs__dfxtp_2
X_4321_ _0620_ u_bits.i_op2\[31\] VSS VSS VCC VCC _1844_ sky130_fd_sc_hs__and2b_1
X_4252_ _1711_ VSS VSS VCC VCC _1800_ sky130_fd_sc_hs__clkbuf_4
X_3203_ _0876_ _0880_ _0825_ VSS VSS VCC VCC _1004_ sky130_fd_sc_hs__mux2_1
X_4183_ _1764_ VSS VSS VCC VCC _0139_ sky130_fd_sc_hs__clkbuf_1
X_3134_ u_muldiv.mul\[25\] _0740_ _0741_ u_muldiv.mul\[57\] _0938_ VSS VSS VCC
+ VCC _0939_ sky130_fd_sc_hs__a221o_1
X_3065_ u_bits.i_op1\[13\] u_bits.i_op1\[12\] _0656_ VSS VSS VCC VCC _0874_
+ sky130_fd_sc_hs__mux2_1
X_3967_ i_rd[1] _1632_ _1636_ o_rd[1] VSS VSS VCC VCC _0051_ sky130_fd_sc_hs__a22o_1
X_5706_ clknet_leaf_30_i_clk _0349_ VSS VSS VCC VCC u_muldiv.quotient_msk\[20\]
+ sky130_fd_sc_hs__dfxtp_1
X_2918_ _0447_ _0727_ _0729_ _0732_ VSS VSS VCC VCC o_result[20] sky130_fd_sc_hs__o211a_2
X_3898_ _1600_ VSS VSS VCC VCC _0018_ sky130_fd_sc_hs__clkbuf_1
X_2849_ _0661_ _0662_ _0663_ VSS VSS VCC VCC _0664_ sky130_fd_sc_hs__mux2_1
X_5637_ clknet_leaf_41_i_clk _0284_ VSS VSS VCC VCC u_muldiv.add_prev\[23\]
+ sky130_fd_sc_hs__dfxtp_1
X_5568_ clknet_leaf_3_i_clk _0215_ VSS VSS VCC VCC u_muldiv.divisor\[49\]
+ sky130_fd_sc_hs__dfxtp_1
X_4519_ _1991_ VSS VSS VCC VCC _0248_ sky130_fd_sc_hs__clkbuf_1
X_5499_ clknet_leaf_43_i_clk _0147_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[17\]
+ sky130_fd_sc_hs__dfxtp_1
X_4870_ _2208_ _2263_ _2264_ _2265_ VSS VSS VCC VCC _2266_ sky130_fd_sc_hs__a31o_1
X_3821_ u_muldiv.mul\[17\] _0717_ _0720_ u_muldiv.mul\[49\] _1540_ VSS VSS VCC
+ VCC _1541_ sky130_fd_sc_hs__a221o_1
X_3752_ _0908_ _1476_ VSS VSS VCC VCC _1477_ sky130_fd_sc_hs__nor2_1
X_3683_ u_muldiv.dividend\[7\] _1326_ _1327_ u_muldiv.o_div\[7\] _1383_ VSS VSS
+ VCC VCC _1413_ sky130_fd_sc_hs__a221o_1
X_2703_ u_bits.i_op1\[12\] u_muldiv.add_prev\[12\] _0450_ VSS VSS VCC VCC
+ _0518_ sky130_fd_sc_hs__mux2_1
X_2634_ _0448_ VSS VSS VCC VCC _0449_ sky130_fd_sc_hs__clkbuf_4
X_5422_ clknet_leaf_48_i_clk _0070_ VSS VSS VCC VCC u_bits.i_op2\[13\] sky130_fd_sc_hs__dfxtp_1
X_5353_ o_add[19] _1214_ VSS VSS VCC VCC _2630_ sky130_fd_sc_hs__and2_1
X_4304_ _1826_ _1827_ VSS VSS VCC VCC _1828_ sky130_fd_sc_hs__nand2_2
X_5284_ u_muldiv.divisor\[0\] _2284_ _2285_ u_muldiv.divisor\[1\] VSS VSS VCC
+ VCC _0391_ sky130_fd_sc_hs__a22o_1
X_4235_ _1791_ VSS VSS VCC VCC _0164_ sky130_fd_sc_hs__clkbuf_1
X_4166_ _1755_ VSS VSS VCC VCC _0131_ sky130_fd_sc_hs__clkbuf_1
X_3117_ _0660_ _0922_ _0664_ _0652_ _0879_ _0923_ VSS VSS VCC VCC _0924_ sky130_fd_sc_hs__mux4_1
X_4097_ u_pc_sel.i_pc_next\[9\] i_pc_next[9] _1712_ VSS VSS VCC VCC _1721_
+ sky130_fd_sc_hs__mux2_1
X_3048_ u_muldiv.mul\[23\] _0717_ _0720_ u_muldiv.mul\[55\] _0856_ VSS VSS VCC
+ VCC _0857_ sky130_fd_sc_hs__a221o_1
X_4999_ u_muldiv.dividend\[6\] _2354_ _2244_ VSS VSS VCC VCC _2355_ sky130_fd_sc_hs__mux2_1
X_4020_ _1487_ _1663_ _1651_ i_op2[13] VSS VSS VCC VCC _1671_ sky130_fd_sc_hs__a22o_1
X_4922_ u_muldiv.quotient_msk\[29\] _2284_ _2283_ u_muldiv.quotient_msk\[30\] VSS
+ VSS VCC VCC _0358_ sky130_fd_sc_hs__a22o_1
X_4853_ u_muldiv.o_div\[24\] _2252_ _2244_ VSS VSS VCC VCC _2253_ sky130_fd_sc_hs__mux2_1
X_4784_ _2170_ u_muldiv.o_div\[11\] _2194_ _2196_ VSS VSS VCC VCC _2197_ sky130_fd_sc_hs__a31o_1
X_3804_ _1524_ _1525_ _0730_ u_pc_sel.i_pc_next\[15\] VSS VSS VCC VCC o_result[15]
+ sky130_fd_sc_hs__a2bb2o_2
X_3735_ _1110_ _1006_ _1458_ _1248_ _1460_ VSS VSS VCC VCC _1461_ sky130_fd_sc_hs__a221o_1
X_5405_ clknet_leaf_51_i_clk _0053_ VSS VSS VCC VCC o_rd[3] sky130_fd_sc_hs__dfxtp_2
X_3666_ _1274_ _1395_ _1396_ _0624_ _1142_ VSS VSS VCC VCC _1397_ sky130_fd_sc_hs__o32a_1
X_3597_ u_muldiv.mul\[2\] _1330_ _1331_ VSS VSS VCC VCC _1332_ sky130_fd_sc_hs__o21ai_1
X_5336_ _1137_ _1585_ VSS VSS VCC VCC _0429_ sky130_fd_sc_hs__nor2_1
X_5267_ _2134_ _2598_ VSS VSS VCC VCC _2599_ sky130_fd_sc_hs__nand2_1
X_4218_ u_wr_mux.i_reg_data2\[26\] i_reg_data2[26] _1778_ VSS VSS VCC VCC
+ _1783_ sky130_fd_sc_hs__mux2_1
X_5198_ u_muldiv.dividend\[24\] _2525_ VSS VSS VCC VCC _2536_ sky130_fd_sc_hs__xor2_1
X_4149_ _1224_ i_funct3[1] _1745_ VSS VSS VCC VCC _1747_ sky130_fd_sc_hs__mux2_1
X_3520_ u_bits.i_op1\[5\] VSS VSS VCC VCC _1257_ sky130_fd_sc_hs__clkbuf_4
X_3451_ u_wr_mux.i_reg_data2\[8\] o_wdata[0] _0718_ VSS VSS VCC VCC _1216_
+ sky130_fd_sc_hs__mux2_1
X_3382_ _1158_ _1161_ VSS VSS VCC VCC _1162_ sky130_fd_sc_hs__xor2_4
X_5121_ _2092_ _2465_ VSS VSS VCC VCC _2466_ sky130_fd_sc_hs__xnor2_1
X_5052_ u_muldiv.dividend\[11\] u_muldiv.dividend\[10\] _2380_ VSS VSS VCC VCC
+ _2403_ sky130_fd_sc_hs__or3_2
X_4003_ u_bits.i_op2\[8\] _1637_ _1651_ i_op2[8] VSS VSS VCC VCC _1659_ sky130_fd_sc_hs__a22o_1
X_4905_ u_muldiv.quotient_msk\[15\] _2280_ _2281_ u_muldiv.quotient_msk\[16\] VSS
+ VSS VCC VCC _0344_ sky130_fd_sc_hs__a22o_1
X_4836_ _2161_ _2238_ u_muldiv.o_div\[21\] VSS VSS VCC VCC _2239_ sky130_fd_sc_hs__a21oi_1
X_4767_ _2167_ _2183_ u_muldiv.o_div\[7\] VSS VSS VCC VCC _2184_ sky130_fd_sc_hs__a21oi_1
X_4698_ _2120_ VSS VSS VCC VCC _2121_ sky130_fd_sc_hs__inv_2
X_3718_ u_bits.i_op2\[10\] VSS VSS VCC VCC _1445_ sky130_fd_sc_hs__clkbuf_4
X_3649_ _1376_ _1257_ _1272_ VSS VSS VCC VCC _1381_ sky130_fd_sc_hs__a21oi_1
X_5319_ _0702_ _1969_ u_bits.i_op2\[31\] VSS VSS VCC VCC _2618_ sky130_fd_sc_hs__a21o_1
X_2951_ _0659_ _0761_ _0762_ _0763_ VSS VSS VCC VCC _0764_ sky130_fd_sc_hs__o22a_1
X_5670_ clknet_leaf_30_i_clk _0313_ VSS VSS VCC VCC u_muldiv.o_div\[16\] sky130_fd_sc_hs__dfxtp_1
X_4621_ u_muldiv.divisor\[12\] u_muldiv.dividend\[12\] VSS VSS VCC VCC _2044_
+ sky130_fd_sc_hs__or2b_1
X_2882_ u_bits.i_op1\[29\] VSS VSS VCC VCC _0697_ sky130_fd_sc_hs__buf_4
X_4552_ _1142_ _2006_ VSS VSS VCC VCC _0266_ sky130_fd_sc_hs__nor2_1
X_4483_ _1972_ VSS VSS VCC VCC _0231_ sky130_fd_sc_hs__clkbuf_1
X_3503_ _1242_ _1243_ VSS VSS VCC VCC o_wsel[0] sky130_fd_sc_hs__nor2_4
X_3434_ i_flush _1203_ VSS VSS VCC VCC _0000_ sky130_fd_sc_hs__nor2_1
X_3365_ _0589_ _1148_ _0603_ VSS VSS VCC VCC _1149_ sky130_fd_sc_hs__a21bo_1
X_5104_ _0654_ _2292_ _2450_ VSS VSS VCC VCC _2451_ sky130_fd_sc_hs__and3_1
X_3296_ _0629_ _1086_ _0955_ VSS VSS VCC VCC _1091_ sky130_fd_sc_hs__a21oi_1
X_5035_ _2295_ _2386_ _1250_ VSS VSS VCC VCC _2388_ sky130_fd_sc_hs__a21oi_1
X_4819_ u_muldiv.o_div\[17\] _2218_ u_muldiv.o_div\[18\] VSS VSS VCC VCC _2225_
+ sky130_fd_sc_hs__o21ai_1
X_5799_ clknet_leaf_34_i_clk _0441_ VSS VSS VCC VCC u_muldiv.mul\[47\] sky130_fd_sc_hs__dfxtp_1
X_3150_ u_mux.i_add_override VSS VSS VCC VCC _0955_ sky130_fd_sc_hs__buf_2
X_3081_ _0730_ _0889_ VSS VSS VCC VCC _0890_ sky130_fd_sc_hs__nor2_1
X_5722_ clknet_leaf_25_i_clk _0365_ VSS VSS VCC VCC u_muldiv.dividend\[6\]
+ sky130_fd_sc_hs__dfxtp_1
X_3983_ _0923_ _1637_ _1638_ i_op2[2] VSS VSS VCC VCC _1645_ sky130_fd_sc_hs__a22o_1
X_2934_ u_mux.i_add_override VSS VSS VCC VCC _0747_ sky130_fd_sc_hs__clkinv_2
X_5653_ clknet_leaf_10_i_clk _0297_ VSS VSS VCC VCC op_cnt\[5\] sky130_fd_sc_hs__dfxtp_1
X_2865_ _0668_ u_bits.i_op1\[0\] _0675_ _0679_ VSS VSS VCC VCC _0680_ sky130_fd_sc_hs__a31o_1
X_4604_ u_muldiv.o_div\[0\] u_muldiv.o_div\[1\] VSS VSS VCC VCC _2027_ sky130_fd_sc_hs__nand2_1
X_5584_ clknet_leaf_38_i_clk _0231_ VSS VSS VCC VCC u_muldiv.mul\[1\] sky130_fd_sc_hs__dfxtp_1
X_4535_ _1999_ VSS VSS VCC VCC _0256_ sky130_fd_sc_hs__clkbuf_1
X_2796_ _0490_ _0491_ VSS VSS VCC VCC _0611_ sky130_fd_sc_hs__or2_1
X_4466_ u_muldiv.divisor\[59\] _1836_ _1946_ u_muldiv.divisor\[60\] _1961_ VSS VSS
+ VCC VCC _0225_ sky130_fd_sc_hs__a221o_1
X_4397_ _1487_ u_bits.i_op2\[14\] _1899_ VSS VSS VCC VCC _1906_ sky130_fd_sc_hs__or3_1
X_3417_ o_add[31] _1185_ _1186_ _1187_ VSS VSS VCC VCC _1188_ sky130_fd_sc_hs__or4_4
X_3348_ _1133_ _1136_ VSS VSS VCC VCC _1137_ sky130_fd_sc_hs__nand2_4
X_3279_ _1015_ _1016_ _1074_ _1047_ VSS VSS VCC VCC _1075_ sky130_fd_sc_hs__a211o_1
X_5018_ _2054_ _2370_ _2288_ VSS VSS VCC VCC _2372_ sky130_fd_sc_hs__a21oi_1
Xclkbuf_0_i_clk i_clk VSS VSS VCC VCC clknet_0_i_clk sky130_fd_sc_hs__clkbuf_16
X_2650_ _0464_ VSS VSS VCC VCC _0465_ sky130_fd_sc_hs__buf_2
X_4320_ _1842_ VSS VSS VCC VCC _1843_ sky130_fd_sc_hs__buf_2
X_4251_ _1799_ VSS VSS VCC VCC _0172_ sky130_fd_sc_hs__clkbuf_1
X_3202_ _0872_ _1002_ _0875_ _0871_ _0879_ _0923_ VSS VSS VCC VCC _1003_ sky130_fd_sc_hs__mux4_1
X_4182_ u_wr_mux.i_reg_data2\[9\] i_reg_data2[9] _1756_ VSS VSS VCC VCC _1764_
+ sky130_fd_sc_hs__mux2_1
X_3133_ u_muldiv.dividend\[25\] _0742_ _0743_ u_muldiv.o_div\[25\] _0744_ VSS VSS
+ VCC VCC _0938_ sky130_fd_sc_hs__a221o_1
X_3064_ _0871_ _0872_ _0696_ VSS VSS VCC VCC _0873_ sky130_fd_sc_hs__mux2_1
X_3966_ i_rd[0] _1632_ _1636_ o_rd[0] VSS VSS VCC VCC _0050_ sky130_fd_sc_hs__a22o_1
X_5705_ clknet_leaf_30_i_clk _0348_ VSS VSS VCC VCC u_muldiv.quotient_msk\[19\]
+ sky130_fd_sc_hs__dfxtp_1
X_2917_ _0731_ VSS VSS VCC VCC _0732_ sky130_fd_sc_hs__buf_2
X_3897_ _1255_ i_op1[2] _1599_ VSS VSS VCC VCC _1600_ sky130_fd_sc_hs__mux2_1
X_5636_ clknet_leaf_42_i_clk _0283_ VSS VSS VCC VCC u_muldiv.add_prev\[22\]
+ sky130_fd_sc_hs__dfxtp_1
X_2848_ _0533_ VSS VSS VCC VCC _0663_ sky130_fd_sc_hs__clkbuf_4
X_2779_ _0592_ _0593_ VSS VSS VCC VCC _0594_ sky130_fd_sc_hs__xnor2_4
X_5567_ clknet_leaf_8_i_clk _0214_ VSS VSS VCC VCC u_muldiv.divisor\[48\]
+ sky130_fd_sc_hs__dfxtp_1
X_4518_ u_muldiv.mul\[18\] u_muldiv.mul\[19\] _1989_ VSS VSS VCC VCC _1991_
+ sky130_fd_sc_hs__mux2_1
X_5498_ clknet_leaf_43_i_clk _0146_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[16\]
+ sky130_fd_sc_hs__dfxtp_1
X_4449_ u_bits.i_op2\[25\] _1947_ VSS VSS VCC VCC _1948_ sky130_fd_sc_hs__nand2_1
X_3820_ u_muldiv.dividend\[17\] _0721_ _0723_ u_muldiv.o_div\[17\] _0724_ VSS VSS
+ VCC VCC _1540_ sky130_fd_sc_hs__a221o_1
X_3751_ _1110_ _1033_ _1473_ _1248_ _1475_ VSS VSS VCC VCC _1476_ sky130_fd_sc_hs__a221o_1
X_2702_ _0457_ _0516_ VSS VSS VCC VCC _0517_ sky130_fd_sc_hs__xnor2_1
X_3682_ _1274_ _1410_ _1411_ _0624_ _1141_ VSS VSS VCC VCC _1412_ sky130_fd_sc_hs__o32a_1
X_2633_ u_mux.i_group_mux VSS VSS VCC VCC _0448_ sky130_fd_sc_hs__buf_2
X_5421_ clknet_leaf_52_i_clk _0069_ VSS VSS VCC VCC u_bits.i_op2\[12\] sky130_fd_sc_hs__dfxtp_4
X_5352_ _2009_ _2628_ VSS VSS VCC VCC _0443_ sky130_fd_sc_hs__nor2_1
X_4303_ u_muldiv.i_on_end VSS VSS VCC VCC _1827_ sky130_fd_sc_hs__clkinv_2
X_5283_ _2164_ _2606_ _2612_ _2613_ VSS VSS VCC VCC _0390_ sky130_fd_sc_hs__a31o_1
X_4234_ csr_data\[0\] i_csr_data[0] _1789_ VSS VSS VCC VCC _1791_ sky130_fd_sc_hs__mux2_1
X_4165_ o_wdata[1] i_reg_data2[1] _1745_ VSS VSS VCC VCC _1755_ sky130_fd_sc_hs__mux2_1
X_3116_ _0825_ VSS VSS VCC VCC _0923_ sky130_fd_sc_hs__clkbuf_4
X_4096_ _1720_ VSS VSS VCC VCC _0096_ sky130_fd_sc_hs__clkbuf_1
X_3047_ u_muldiv.dividend\[23\] _0633_ _0722_ u_muldiv.o_div\[23\] _0724_ VSS VSS
+ VCC VCC _0856_ sky130_fd_sc_hs__a221o_1
X_4998_ _1208_ _2345_ _2346_ _2353_ VSS VSS VCC VCC _2354_ sky130_fd_sc_hs__a31o_1
X_3949_ _0996_ i_op1[27] _1621_ VSS VSS VCC VCC _1627_ sky130_fd_sc_hs__mux2_1
X_5619_ clknet_leaf_45_i_clk _0266_ VSS VSS VCC VCC u_muldiv.add_prev\[5\]
+ sky130_fd_sc_hs__dfxtp_1
Xclkbuf_leaf_16_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_16_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4921_ u_muldiv.quotient_msk\[28\] _2284_ _2283_ u_muldiv.quotient_msk\[29\] VSS
+ VSS VCC VCC _0357_ sky130_fd_sc_hs__a22o_1
X_4852_ _2208_ _2249_ _2250_ _2251_ VSS VSS VCC VCC _2252_ sky130_fd_sc_hs__a31o_1
X_3803_ _1333_ csr_data\[15\] _0731_ VSS VSS VCC VCC _1525_ sky130_fd_sc_hs__o21ai_1
X_4783_ _1880_ VSS VSS VCC VCC _2196_ sky130_fd_sc_hs__clkbuf_4
X_3734_ u_bits.i_op2\[11\] _1251_ _0926_ _1459_ VSS VSS VCC VCC _1460_ sky130_fd_sc_hs__o22a_1
X_3665_ u_bits.i_op2\[6\] _0786_ _1272_ VSS VSS VCC VCC _1396_ sky130_fd_sc_hs__a21oi_1
X_5404_ clknet_leaf_51_i_clk _0052_ VSS VSS VCC VCC o_rd[2] sky130_fd_sc_hs__dfxtp_2
X_3596_ _0453_ VSS VSS VCC VCC _1331_ sky130_fd_sc_hs__buf_2
X_5335_ _1128_ _1585_ VSS VSS VCC VCC _0428_ sky130_fd_sc_hs__nor2_1
X_5266_ _2030_ _2131_ _2132_ _2133_ VSS VSS VCC VCC _2598_ sky130_fd_sc_hs__a31o_1
X_4217_ _1782_ VSS VSS VCC VCC _0155_ sky130_fd_sc_hs__clkbuf_1
X_5197_ _2535_ VSS VSS VCC VCC _0382_ sky130_fd_sc_hs__clkbuf_1
X_4148_ _1746_ VSS VSS VCC VCC _0122_ sky130_fd_sc_hs__clkbuf_1
X_4079_ _1594_ VSS VSS VCC VCC _1711_ sky130_fd_sc_hs__buf_4
X_3450_ _1215_ VSS VSS VCC VCC _0003_ sky130_fd_sc_hs__clkbuf_1
X_3381_ _1159_ _1160_ _0507_ VSS VSS VCC VCC _1161_ sky130_fd_sc_hs__a21bo_1
X_5120_ _2458_ _2089_ _2087_ VSS VSS VCC VCC _2465_ sky130_fd_sc_hs__o21a_1
X_5051_ _2402_ VSS VSS VCC VCC _0369_ sky130_fd_sc_hs__clkbuf_1
X_4002_ u_bits.i_op2\[9\] _1406_ _1657_ VSS VSS VCC VCC _1658_ sky130_fd_sc_hs__mux2_1
X_4904_ u_muldiv.quotient_msk\[14\] _2280_ _2281_ u_muldiv.quotient_msk\[15\] VSS
+ VSS VCC VCC _0343_ sky130_fd_sc_hs__a22o_1
X_4835_ u_muldiv.quotient_msk\[21\] _2233_ _2229_ VSS VSS VCC VCC _2238_ sky130_fd_sc_hs__mux2_1
X_4766_ u_muldiv.quotient_msk\[7\] _2179_ _2156_ VSS VSS VCC VCC _2183_ sky130_fd_sc_hs__mux2_1
X_3717_ _1443_ _1315_ _0970_ _0824_ _0670_ _0643_ VSS VSS VCC VCC _1444_ sky130_fd_sc_hs__mux4_1
X_4697_ u_muldiv.dividend\[23\] u_muldiv.divisor\[23\] VSS VSS VCC VCC _2120_
+ sky130_fd_sc_hs__and2b_1
X_3648_ _1249_ _1375_ _1379_ VSS VSS VCC VCC _1380_ sky130_fd_sc_hs__a21oi_1
X_3579_ _0645_ _0646_ _0630_ _0768_ _0658_ _0659_ VSS VSS VCC VCC _1314_ sky130_fd_sc_hs__mux4_1
X_5318_ u_muldiv.divisor\[30\] _1838_ _1843_ u_muldiv.divisor\[31\] VSS VSS VCC
+ VCC _0421_ sky130_fd_sc_hs__a22o_1
X_5249_ _2582_ VSS VSS VCC VCC _0387_ sky130_fd_sc_hs__clkbuf_1
X_2950_ _0657_ _0702_ VSS VSS VCC VCC _0763_ sky130_fd_sc_hs__and2b_1
X_2881_ u_bits.i_op2\[2\] VSS VSS VCC VCC _0696_ sky130_fd_sc_hs__buf_4
X_4620_ u_muldiv.dividend\[13\] u_muldiv.divisor\[13\] VSS VSS VCC VCC _2043_
+ sky130_fd_sc_hs__and2b_1
X_4551_ _1135_ _2006_ VSS VSS VCC VCC _0265_ sky130_fd_sc_hs__nor2_1
X_4482_ u_muldiv.mul\[1\] u_muldiv.mul\[2\] _1584_ VSS VSS VCC VCC _1972_
+ sky130_fd_sc_hs__mux2_1
X_3502_ _1233_ o_add[0] VSS VSS VCC VCC _1243_ sky130_fd_sc_hs__and2_1
X_3433_ u_muldiv.i_on_wait _1202_ VSS VSS VCC VCC _1203_ sky130_fd_sc_hs__nand2_1
X_3364_ _0594_ _1143_ _0605_ VSS VSS VCC VCC _1148_ sky130_fd_sc_hs__o21ai_2
X_5103_ u_bits.i_op1\[13\] u_bits.i_op1\[14\] _2428_ VSS VSS VCC VCC _2450_
+ sky130_fd_sc_hs__or3_2
X_3295_ _0628_ _1082_ _1089_ VSS VSS VCC VCC _1090_ sky130_fd_sc_hs__or3_2
X_5034_ _1250_ _2385_ _2386_ VSS VSS VCC VCC _2387_ sky130_fd_sc_hs__and3_1
X_4818_ _2181_ _2222_ _2224_ VSS VSS VCC VCC _0314_ sky130_fd_sc_hs__a21oi_1
X_5798_ clknet_leaf_39_i_clk _0440_ VSS VSS VCC VCC u_muldiv.mul\[46\] sky130_fd_sc_hs__dfxtp_1
X_4749_ _2164_ _2166_ _2169_ VSS VSS VCC VCC _0300_ sky130_fd_sc_hs__a21oi_1
X_3080_ _0857_ _0888_ _0446_ VSS VSS VCC VCC _0889_ sky130_fd_sc_hs__a21oi_2
X_3982_ _0909_ _1112_ _1639_ VSS VSS VCC VCC _1644_ sky130_fd_sc_hs__mux2_1
X_5721_ clknet_leaf_25_i_clk _0364_ VSS VSS VCC VCC u_muldiv.dividend\[5\]
+ sky130_fd_sc_hs__dfxtp_1
X_2933_ u_muldiv.mul\[21\] _0740_ _0741_ u_muldiv.mul\[53\] _0745_ VSS VSS VCC
+ VCC _0746_ sky130_fd_sc_hs__a221o_1
X_5652_ clknet_leaf_10_i_clk _0296_ VSS VSS VCC VCC op_cnt\[4\] sky130_fd_sc_hs__dfxtp_1
X_2864_ u_bits.i_op2\[2\] _0678_ VSS VSS VCC VCC _0679_ sky130_fd_sc_hs__and2b_1
X_4603_ u_muldiv.o_div\[0\] u_muldiv.o_div\[1\] VSS VSS VCC VCC _2026_ sky130_fd_sc_hs__or2_1
X_5583_ clknet_leaf_35_i_clk _0230_ VSS VSS VCC VCC u_muldiv.mul\[0\] sky130_fd_sc_hs__dfxtp_1
X_2795_ _0488_ _0609_ VSS VSS VCC VCC _0610_ sky130_fd_sc_hs__nand2_1
X_4534_ u_muldiv.mul\[26\] u_muldiv.mul\[27\] _1989_ VSS VSS VCC VCC _1999_
+ sky130_fd_sc_hs__mux2_1
X_4465_ _1959_ _1960_ VSS VSS VCC VCC _1961_ sky130_fd_sc_hs__nor2_1
X_3416_ o_add[29] o_add[30] VSS VSS VCC VCC _1187_ sky130_fd_sc_hs__or2_1
X_4396_ u_muldiv.divisor\[45\] _1867_ _1887_ u_muldiv.divisor\[46\] _1905_ VSS VSS
+ VCC VCC _0211_ sky130_fd_sc_hs__a221o_1
X_3347_ _1131_ _1132_ VSS VSS VCC VCC _1136_ sky130_fd_sc_hs__or2_1
X_5017_ _2054_ _2370_ VSS VSS VCC VCC _2371_ sky130_fd_sc_hs__or2_1
X_3278_ _1023_ VSS VSS VCC VCC _1074_ sky130_fd_sc_hs__inv_2
X_4250_ csr_data\[8\] i_csr_data[8] _1789_ VSS VSS VCC VCC _1799_ sky130_fd_sc_hs__mux2_1
X_4181_ _1763_ VSS VSS VCC VCC _0138_ sky130_fd_sc_hs__clkbuf_1
X_3201_ _1001_ _0944_ _0774_ VSS VSS VCC VCC _1002_ sky130_fd_sc_hs__mux2_1
X_3132_ _0936_ _0937_ VSS VSS VCC VCC o_add[25] sky130_fd_sc_hs__xnor2_4
X_3063_ _0773_ _0781_ _0533_ VSS VSS VCC VCC _0872_ sky130_fd_sc_hs__mux2_1
X_3965_ i_reg_write _1632_ _1636_ o_reg_write VSS VSS VCC VCC _0049_ sky130_fd_sc_hs__a22o_1
X_5704_ clknet_leaf_30_i_clk _0347_ VSS VSS VCC VCC u_muldiv.quotient_msk\[18\]
+ sky130_fd_sc_hs__dfxtp_1
X_2916_ _0730_ VSS VSS VCC VCC _0731_ sky130_fd_sc_hs__inv_2
X_3896_ _1595_ VSS VSS VCC VCC _1599_ sky130_fd_sc_hs__clkbuf_4
X_2847_ u_bits.i_op1\[10\] u_bits.i_op1\[9\] _0649_ VSS VSS VCC VCC _0662_
+ sky130_fd_sc_hs__mux2_1
X_5635_ clknet_leaf_41_i_clk _0282_ VSS VSS VCC VCC u_muldiv.add_prev\[21\]
+ sky130_fd_sc_hs__dfxtp_1
X_2778_ u_bits.i_op1\[9\] u_muldiv.add_prev\[9\] _0450_ VSS VSS VCC VCC _0593_
+ sky130_fd_sc_hs__mux2_2
X_5566_ clknet_leaf_8_i_clk _0213_ VSS VSS VCC VCC u_muldiv.divisor\[47\]
+ sky130_fd_sc_hs__dfxtp_1
X_4517_ _1990_ VSS VSS VCC VCC _0247_ sky130_fd_sc_hs__clkbuf_1
X_5497_ clknet_leaf_43_i_clk _0145_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[15\]
+ sky130_fd_sc_hs__dfxtp_1
X_4448_ _0905_ _1942_ _1846_ VSS VSS VCC VCC _1947_ sky130_fd_sc_hs__o21ai_1
X_4379_ _1445_ _1888_ _1846_ VSS VSS VCC VCC _1892_ sky130_fd_sc_hs__o21a_1
X_3750_ u_bits.i_op2\[12\] _0777_ _0926_ _1474_ VSS VSS VCC VCC _1475_ sky130_fd_sc_hs__o22a_1
X_2701_ _0460_ u_bits.i_op2\[12\] u_bits.i_op1\[12\] _0464_ VSS VSS VCC VCC
+ _0516_ sky130_fd_sc_hs__a22o_1
X_3681_ _1406_ _1258_ _1272_ VSS VSS VCC VCC _1411_ sky130_fd_sc_hs__a21oi_1
X_2632_ _0446_ VSS VSS VCC VCC _0447_ sky130_fd_sc_hs__clkbuf_4
X_5420_ clknet_leaf_52_i_clk _0068_ VSS VSS VCC VCC u_bits.i_op2\[11\] sky130_fd_sc_hs__dfxtp_4
X_5351_ _1176_ _2628_ VSS VSS VCC VCC _0442_ sky130_fd_sc_hs__nor2_1
X_4302_ u_muldiv.on_wait VSS VSS VCC VCC _1826_ sky130_fd_sc_hs__clkbuf_4
X_5282_ u_muldiv.dividend\[31\] _2157_ VSS VSS VCC VCC _2613_ sky130_fd_sc_hs__and2_1
X_4233_ i_to_trap _1638_ _1635_ o_to_trap VSS VSS VCC VCC _0163_ sky130_fd_sc_hs__a22o_1
X_4164_ _1754_ VSS VSS VCC VCC _0130_ sky130_fd_sc_hs__clkbuf_1
X_4095_ u_pc_sel.i_pc_next\[8\] i_pc_next[8] _1712_ VSS VSS VCC VCC _1720_
+ sky130_fd_sc_hs__mux2_1
X_3115_ _0904_ _0692_ _0691_ _0768_ _0658_ _0659_ VSS VSS VCC VCC _0922_ sky130_fd_sc_hs__mux4_1
X_3046_ _0855_ VSS VSS VCC VCC o_add[23] sky130_fd_sc_hs__inv_2
X_4997_ _1207_ _2352_ VSS VSS VCC VCC _2353_ sky130_fd_sc_hs__nor2_1
X_3948_ _1626_ VSS VSS VCC VCC _0042_ sky130_fd_sc_hs__clkbuf_1
X_3879_ o_add[29] _1579_ VSS VSS VCC VCC _1588_ sky130_fd_sc_hs__and2_1
X_5618_ clknet_leaf_45_i_clk _0265_ VSS VSS VCC VCC u_muldiv.add_prev\[4\]
+ sky130_fd_sc_hs__dfxtp_1
X_5549_ clknet_leaf_6_i_clk mul_op2_signed_next VSS VSS VCC VCC u_muldiv.i_op2_signed
+ sky130_fd_sc_hs__dfxtp_1
X_4920_ u_muldiv.quotient_msk\[27\] _2284_ _2283_ u_muldiv.quotient_msk\[28\] VSS
+ VSS VCC VCC _0356_ sky130_fd_sc_hs__a22o_1
X_4851_ u_muldiv.quotient_msk\[24\] u_muldiv.o_div\[24\] _1840_ VSS VSS VCC
+ VCC _2251_ sky130_fd_sc_hs__o21a_1
X_3802_ _1331_ _1520_ _1522_ _1523_ _0728_ VSS VSS VCC VCC _1524_ sky130_fd_sc_hs__o221a_1
X_4782_ u_muldiv.o_div\[10\] _2171_ _2195_ _2164_ VSS VSS VCC VCC _0307_ sky130_fd_sc_hs__a22o_1
X_3733_ u_bits.i_op2\[11\] _1251_ _1267_ VSS VSS VCC VCC _1459_ sky130_fd_sc_hs__a21oi_1
X_3664_ _1249_ _1391_ _1394_ VSS VSS VCC VCC _1395_ sky130_fd_sc_hs__a21oi_1
X_5403_ clknet_leaf_51_i_clk _0051_ VSS VSS VCC VCC o_rd[1] sky130_fd_sc_hs__dfxtp_2
X_3595_ _0748_ VSS VSS VCC VCC _1330_ sky130_fd_sc_hs__buf_2
X_5334_ _1130_ _1585_ VSS VSS VCC VCC _0427_ sky130_fd_sc_hs__nor2_1
X_5265_ _2375_ _2135_ VSS VSS VCC VCC _2597_ sky130_fd_sc_hs__nor2_1
X_5196_ u_muldiv.dividend\[23\] _2534_ _2485_ VSS VSS VCC VCC _2535_ sky130_fd_sc_hs__mux2_1
X_4216_ u_wr_mux.i_reg_data2\[25\] i_reg_data2[25] _1778_ VSS VSS VCC VCC
+ _1782_ sky130_fd_sc_hs__mux2_1
X_4147_ _0620_ i_funct3[0] _1745_ VSS VSS VCC VCC _1746_ sky130_fd_sc_hs__mux2_1
X_4078_ u_bits.i_op2\[30\] _1639_ _1635_ _1710_ VSS VSS VCC VCC _0088_ sky130_fd_sc_hs__a31o_1
X_3029_ _0677_ _0839_ _0779_ VSS VSS VCC VCC _0840_ sky130_fd_sc_hs__mux2_1
X_3380_ _0577_ _1153_ _0521_ VSS VSS VCC VCC _1160_ sky130_fd_sc_hs__o21ai_2
X_5050_ u_muldiv.dividend\[10\] _2401_ _2378_ VSS VSS VCC VCC _2402_ sky130_fd_sc_hs__mux2_1
X_4001_ _1198_ VSS VSS VCC VCC _1657_ sky130_fd_sc_hs__clkbuf_4
X_4903_ u_muldiv.quotient_msk\[13\] _2280_ _2281_ u_muldiv.quotient_msk\[14\] VSS
+ VSS VCC VCC _0342_ sky130_fd_sc_hs__a22o_1
X_4834_ u_muldiv.o_div\[21\] _2170_ _2233_ _2196_ VSS VSS VCC VCC _2237_ sky130_fd_sc_hs__a31o_1
X_4765_ _2165_ u_muldiv.o_div\[7\] _2179_ _1913_ VSS VSS VCC VCC _2182_ sky130_fd_sc_hs__a31o_1
X_3716_ _1306_ _1309_ _0760_ VSS VSS VCC VCC _1443_ sky130_fd_sc_hs__mux2_1
X_4696_ _2112_ _2118_ VSS VSS VCC VCC _2119_ sky130_fd_sc_hs__nor2_1
Xclkbuf_leaf_15_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_15_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3647_ _1265_ _0797_ _1378_ _0634_ VSS VSS VCC VCC _1379_ sky130_fd_sc_hs__o211ai_1
X_3578_ _1306_ _1309_ _1311_ _1312_ _0789_ _0674_ VSS VSS VCC VCC _1313_ sky130_fd_sc_hs__mux4_1
X_5317_ u_muldiv.divisor\[29\] _1838_ _1843_ u_muldiv.divisor\[30\] VSS VSS VCC
+ VCC _0420_ sky130_fd_sc_hs__a22o_1
X_5248_ u_muldiv.dividend\[28\] _2581_ _2485_ VSS VSS VCC VCC _2582_ sky130_fd_sc_hs__mux2_1
X_5179_ _0768_ _2511_ _2385_ VSS VSS VCC VCC _2519_ sky130_fd_sc_hs__o21ai_1
X_2880_ _0669_ _0690_ _0694_ VSS VSS VCC VCC _0695_ sky130_fd_sc_hs__a21oi_1
X_4550_ _1137_ _2006_ VSS VSS VCC VCC _0264_ sky130_fd_sc_hs__nor2_1
X_4481_ _1971_ VSS VSS VCC VCC _0230_ sky130_fd_sc_hs__clkbuf_1
X_3501_ _0619_ o_add[1] VSS VSS VCC VCC _1242_ sky130_fd_sc_hs__and2b_1
X_3432_ _1199_ _1201_ op_cnt\[0\] VSS VSS VCC VCC _1202_ sky130_fd_sc_hs__a21oi_1
X_3363_ _1147_ VSS VSS VCC VCC o_add[8] sky130_fd_sc_hs__inv_2
X_5102_ _2447_ _2448_ VSS VSS VCC VCC _2449_ sky130_fd_sc_hs__xnor2_1
X_3294_ _0925_ _1084_ _1085_ _0914_ _1088_ VSS VSS VCC VCC _1089_ sky130_fd_sc_hs__a221o_1
X_5033_ u_bits.i_op1\[7\] u_bits.i_op1\[8\] _2363_ VSS VSS VCC VCC _2386_
+ sky130_fd_sc_hs__or3_2
X_4817_ _2161_ _2223_ u_muldiv.o_div\[17\] VSS VSS VCC VCC _2224_ sky130_fd_sc_hs__a21oi_1
X_5797_ clknet_leaf_39_i_clk _0439_ VSS VSS VCC VCC u_muldiv.mul\[45\] sky130_fd_sc_hs__dfxtp_1
X_4748_ _2167_ _2168_ u_muldiv.o_div\[3\] VSS VSS VCC VCC _2169_ sky130_fd_sc_hs__a21oi_1
X_4679_ _2036_ _2038_ _2098_ _2101_ VSS VSS VCC VCC _2102_ sky130_fd_sc_hs__a31o_1
X_3981_ _1641_ _1642_ _1643_ VSS VSS VCC VCC _0058_ sky130_fd_sc_hs__a21o_1
X_2932_ u_muldiv.dividend\[21\] _0742_ _0743_ u_muldiv.o_div\[21\] _0744_ VSS VSS
+ VCC VCC _0745_ sky130_fd_sc_hs__a221o_1
X_5720_ clknet_leaf_25_i_clk _0363_ VSS VSS VCC VCC u_muldiv.dividend\[4\]
+ sky130_fd_sc_hs__dfxtp_1
X_5651_ clknet_leaf_10_i_clk _0295_ VSS VSS VCC VCC op_cnt\[3\] sky130_fd_sc_hs__dfxtp_1
X_2863_ _0676_ _0677_ _0533_ VSS VSS VCC VCC _0678_ sky130_fd_sc_hs__mux2_1
X_4602_ op_cnt\[5\] _2023_ _2025_ VSS VSS VCC VCC _0297_ sky130_fd_sc_hs__o21a_1
X_5582_ clknet_leaf_36_i_clk _0229_ VSS VSS VCC VCC u_muldiv.quotient_msk\[31\]
+ sky130_fd_sc_hs__dfxtp_1
X_2794_ _0493_ VSS VSS VCC VCC _0609_ sky130_fd_sc_hs__inv_2
X_4533_ _1998_ VSS VSS VCC VCC _0255_ sky130_fd_sc_hs__clkbuf_1
X_4464_ u_bits.i_op2\[28\] _1852_ _1958_ _1856_ VSS VSS VCC VCC _1960_ sky130_fd_sc_hs__a31o_1
X_3415_ _0993_ _1024_ VSS VSS VCC VCC _1186_ sky130_fd_sc_hs__nand2_1
X_4395_ _1832_ _1904_ VSS VSS VCC VCC _1905_ sky130_fd_sc_hs__nor2_1
X_3346_ _1135_ VSS VSS VCC VCC o_add[5] sky130_fd_sc_hs__inv_2
X_5016_ _2055_ _2075_ VSS VSS VCC VCC _2370_ sky130_fd_sc_hs__or2_1
X_3277_ _1045_ VSS VSS VCC VCC _1073_ sky130_fd_sc_hs__inv_2
X_4180_ u_wr_mux.i_reg_data2\[8\] i_reg_data2[8] _1756_ VSS VSS VCC VCC _1763_
+ sky130_fd_sc_hs__mux2_1
X_3200_ u_bits.i_op1\[27\] _0689_ _0778_ VSS VSS VCC VCC _1001_ sky130_fd_sc_hs__mux2_1
X_3131_ _0898_ _0899_ _0901_ VSS VSS VCC VCC _0937_ sky130_fd_sc_hs__a21bo_1
X_3062_ _0870_ _0772_ _0533_ VSS VSS VCC VCC _0871_ sky130_fd_sc_hs__mux2_1
X_3964_ i_store _1632_ _1636_ o_store VSS VSS VCC VCC _0048_ sky130_fd_sc_hs__a22o_1
X_5703_ clknet_leaf_30_i_clk _0346_ VSS VSS VCC VCC u_muldiv.quotient_msk\[17\]
+ sky130_fd_sc_hs__dfxtp_1
X_2915_ o_res_src[1] VSS VSS VCC VCC _0730_ sky130_fd_sc_hs__buf_2
X_3895_ _1598_ VSS VSS VCC VCC _0017_ sky130_fd_sc_hs__clkbuf_1
X_2846_ u_bits.i_op1\[12\] u_bits.i_op1\[11\] _0657_ VSS VSS VCC VCC _0661_
+ sky130_fd_sc_hs__mux2_1
X_5634_ clknet_leaf_41_i_clk _0281_ VSS VSS VCC VCC u_muldiv.add_prev\[20\]
+ sky130_fd_sc_hs__dfxtp_1
X_2777_ _0457_ _0591_ VSS VSS VCC VCC _0592_ sky130_fd_sc_hs__xnor2_4
X_5565_ clknet_leaf_8_i_clk _0212_ VSS VSS VCC VCC u_muldiv.divisor\[46\]
+ sky130_fd_sc_hs__dfxtp_1
X_4516_ u_muldiv.mul\[17\] u_muldiv.mul\[18\] _1989_ VSS VSS VCC VCC _1990_
+ sky130_fd_sc_hs__mux2_1
X_5496_ clknet_leaf_43_i_clk _0144_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[14\]
+ sky130_fd_sc_hs__dfxtp_1
X_4447_ _1841_ VSS VSS VCC VCC _1946_ sky130_fd_sc_hs__buf_4
X_4378_ u_muldiv.divisor\[41\] _1867_ _1887_ u_muldiv.divisor\[42\] _1891_ VSS VSS
+ VCC VCC _0207_ sky130_fd_sc_hs__a221o_1
X_3329_ _0749_ o_add[31] _1120_ _1121_ _0453_ VSS VSS VCC VCC _1122_ sky130_fd_sc_hs__a221o_1
X_2700_ _0513_ _0514_ VSS VSS VCC VCC _0515_ sky130_fd_sc_hs__nor2_1
X_3680_ _1249_ _1405_ _1409_ VSS VSS VCC VCC _1410_ sky130_fd_sc_hs__a21oi_1
X_2631_ csr_read VSS VSS VCC VCC _0446_ sky130_fd_sc_hs__buf_4
X_5350_ _2629_ VSS VSS VCC VCC _0441_ sky130_fd_sc_hs__clkbuf_1
X_5281_ _2303_ _2609_ _2611_ _2165_ VSS VSS VCC VCC _2612_ sky130_fd_sc_hs__a211o_1
X_4301_ i_inst_branch i_funct3[0] _1632_ _1825_ VSS VSS VCC VCC _0196_ sky130_fd_sc_hs__a31o_1
X_4232_ _1790_ VSS VSS VCC VCC _0162_ sky130_fd_sc_hs__clkbuf_1
X_4163_ o_wdata[0] i_reg_data2[0] _1745_ VSS VSS VCC VCC _1754_ sky130_fd_sc_hs__mux2_1
X_3114_ _0916_ _0918_ _0919_ _0920_ VSS VSS VCC VCC _0921_ sky130_fd_sc_hs__a2bb2o_1
X_4094_ _1719_ VSS VSS VCC VCC _0095_ sky130_fd_sc_hs__clkbuf_1
X_3045_ _0853_ _0854_ VSS VSS VCC VCC _0855_ sky130_fd_sc_hs__xnor2_2
X_4996_ _2347_ _2349_ _2351_ _1826_ VSS VSS VCC VCC _2352_ sky130_fd_sc_hs__o22a_1
X_3947_ _0689_ i_op1[26] _1621_ VSS VSS VCC VCC _1626_ sky130_fd_sc_hs__mux2_1
X_3878_ _1024_ _1585_ VSS VSS VCC VCC _0011_ sky130_fd_sc_hs__nor2_1
X_5617_ clknet_leaf_45_i_clk _0264_ VSS VSS VCC VCC u_muldiv.add_prev\[3\]
+ sky130_fd_sc_hs__dfxtp_1
X_2829_ _0643_ VSS VSS VCC VCC _0644_ sky130_fd_sc_hs__clkbuf_4
X_5548_ clknet_leaf_5_i_clk _0196_ VSS VSS VCC VCC u_adder.i_cmp_inverse sky130_fd_sc_hs__dfxtp_1
X_5479_ clknet_leaf_6_i_clk _0127_ VSS VSS VCC VCC alu_ctrl\[2\] sky130_fd_sc_hs__dfxtp_1
X_4850_ u_muldiv.o_div\[23\] u_muldiv.o_div\[24\] _2241_ VSS VSS VCC VCC _2250_
+ sky130_fd_sc_hs__or3_2
X_3801_ u_muldiv.mul\[15\] _0748_ _1400_ VSS VSS VCC VCC _1523_ sky130_fd_sc_hs__o21ai_1
X_4781_ _2165_ _2193_ _2194_ _1842_ u_muldiv.quotient_msk\[10\] VSS VSS VCC
+ VCC _2195_ sky130_fd_sc_hs__a32o_1
X_3732_ _1457_ _1344_ _0998_ _0824_ _0707_ _0643_ VSS VSS VCC VCC _1458_ sky130_fd_sc_hs__mux4_1
X_3663_ _0674_ _1110_ _0841_ _1393_ _0858_ VSS VSS VCC VCC _1394_ sky130_fd_sc_hs__a311o_1
X_5402_ clknet_leaf_51_i_clk _0050_ VSS VSS VCC VCC o_rd[0] sky130_fd_sc_hs__dfxtp_2
X_3594_ u_muldiv.mul\[34\] _1325_ _1328_ VSS VSS VCC VCC _1329_ sky130_fd_sc_hs__a21oi_1
X_5333_ _2627_ VSS VSS VCC VCC _0426_ sky130_fd_sc_hs__clkbuf_1
X_5264_ _0699_ _2362_ _2594_ VSS VSS VCC VCC _2596_ sky130_fd_sc_hs__nand3_1
X_5195_ _1208_ _2525_ _2526_ _2533_ VSS VSS VCC VCC _2534_ sky130_fd_sc_hs__a31o_1
X_4215_ _1781_ VSS VSS VCC VCC _0154_ sky130_fd_sc_hs__clkbuf_1
X_4146_ _1711_ VSS VSS VCC VCC _1745_ sky130_fd_sc_hs__buf_4
X_4077_ u_bits.i_op2\[31\] _1634_ _1596_ i_op2[31] VSS VSS VCC VCC _1710_
+ sky130_fd_sc_hs__a22o_1
X_3028_ _0658_ u_bits.i_op1\[0\] VSS VSS VCC VCC _0839_ sky130_fd_sc_hs__and2b_1
X_4979_ u_muldiv.dividend\[5\] u_muldiv.dividend\[4\] _2315_ VSS VSS VCC VCC
+ _2336_ sky130_fd_sc_hs__or3_1
X_4000_ _1641_ _1655_ _1656_ VSS VSS VCC VCC _0064_ sky130_fd_sc_hs__a21o_1
X_4902_ u_muldiv.quotient_msk\[12\] _2280_ _2281_ u_muldiv.quotient_msk\[13\] VSS
+ VSS VCC VCC _0341_ sky130_fd_sc_hs__a22o_1
X_4833_ _2236_ VSS VSS VCC VCC _0317_ sky130_fd_sc_hs__clkbuf_1
X_4764_ _2154_ VSS VSS VCC VCC _2181_ sky130_fd_sc_hs__buf_2
X_3715_ _1441_ _1442_ _1336_ u_pc_sel.i_pc_next\[9\] VSS VSS VCC VCC o_result[9]
+ sky130_fd_sc_hs__a2bb2o_2
X_4695_ _2113_ _2117_ VSS VSS VCC VCC _2118_ sky130_fd_sc_hs__nand2_1
X_3646_ _1376_ _1257_ _1293_ _1377_ VSS VSS VCC VCC _1378_ sky130_fd_sc_hs__a2bb2o_1
X_3577_ _0786_ _1258_ _0785_ _1250_ _0651_ _0774_ VSS VSS VCC VCC _1312_ sky130_fd_sc_hs__mux4_1
X_5316_ u_muldiv.divisor\[28\] _1838_ _2617_ u_muldiv.divisor\[29\] VSS VSS VCC
+ VCC _0419_ sky130_fd_sc_hs__a22o_1
X_5247_ _2575_ _2579_ _1877_ _2580_ VSS VSS VCC VCC _2581_ sky130_fd_sc_hs__o2bb2a_1
X_5178_ _2104_ _2035_ _2102_ _1839_ VSS VSS VCC VCC _2518_ sky130_fd_sc_hs__a31o_1
X_4129_ _1736_ VSS VSS VCC VCC _0113_ sky130_fd_sc_hs__clkbuf_1
X_3500_ _1192_ u_wr_mux.i_reg_data2\[31\] _1241_ VSS VSS VCC VCC o_wdata[31]
+ sky130_fd_sc_hs__a21o_2
X_4480_ u_muldiv.mul\[0\] u_muldiv.mul\[1\] _1584_ VSS VSS VCC VCC _1971_
+ sky130_fd_sc_hs__mux2_1
X_3431_ _1198_ op_cnt\[5\] _1200_ op_cnt\[4\] VSS VSS VCC VCC _1201_ sky130_fd_sc_hs__or4b_1
X_3362_ _1143_ _1146_ VSS VSS VCC VCC _1147_ sky130_fd_sc_hs__nand2_2
X_5101_ _2039_ _2082_ VSS VSS VCC VCC _2448_ sky130_fd_sc_hs__and2b_1
X_3293_ _0699_ u_bits.i_op2\[30\] _0636_ _1087_ VSS VSS VCC VCC _1088_ sky130_fd_sc_hs__o22a_1
X_5032_ _2292_ VSS VSS VCC VCC _2385_ sky130_fd_sc_hs__buf_2
X_4816_ u_muldiv.quotient_msk\[17\] _2218_ _2156_ VSS VSS VCC VCC _2223_ sky130_fd_sc_hs__mux2_1
X_5796_ clknet_leaf_34_i_clk _0438_ VSS VSS VCC VCC u_muldiv.mul\[44\] sky130_fd_sc_hs__dfxtp_1
X_4747_ u_muldiv.quotient_msk\[3\] _2158_ _2156_ VSS VSS VCC VCC _2168_ sky130_fd_sc_hs__mux2_1
X_4678_ _2034_ _2100_ _2032_ VSS VSS VCC VCC _2101_ sky130_fd_sc_hs__or3b_1
X_3629_ _0751_ _0708_ _1361_ _0710_ VSS VSS VCC VCC _1362_ sky130_fd_sc_hs__a211o_1
Xclkbuf_leaf_14_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_14_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3980_ _1112_ _1637_ _1638_ i_op2[1] VSS VSS VCC VCC _1643_ sky130_fd_sc_hs__a22o_1
X_2931_ _0724_ VSS VSS VCC VCC _0744_ sky130_fd_sc_hs__clkbuf_4
X_5650_ clknet_leaf_11_i_clk _0294_ VSS VSS VCC VCC op_cnt\[2\] sky130_fd_sc_hs__dfxtp_1
X_4601_ op_cnt\[5\] _2023_ _1204_ VSS VSS VCC VCC _2025_ sky130_fd_sc_hs__a21oi_1
X_2862_ u_bits.i_op1\[2\] u_bits.i_op1\[1\] _0656_ VSS VSS VCC VCC _0677_
+ sky130_fd_sc_hs__mux2_1
Xclkbuf_leaf_29_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_29_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_2793_ _0579_ _0607_ VSS VSS VCC VCC _0608_ sky130_fd_sc_hs__or2_1
X_5581_ clknet_leaf_3_i_clk _0228_ VSS VSS VCC VCC u_muldiv.divisor\[62\]
+ sky130_fd_sc_hs__dfxtp_1
X_4532_ u_muldiv.mul\[25\] u_muldiv.mul\[26\] _1989_ VSS VSS VCC VCC _1998_
+ sky130_fd_sc_hs__mux2_1
X_4463_ _1868_ _1958_ u_bits.i_op2\[28\] VSS VSS VCC VCC _1959_ sky130_fd_sc_hs__a21oi_1
X_3414_ o_add[25] o_add[26] _1183_ _1184_ VSS VSS VCC VCC _1185_ sky130_fd_sc_hs__or4_1
X_4394_ u_bits.i_op2\[14\] _1903_ VSS VSS VCC VCC _1904_ sky130_fd_sc_hs__xnor2_1
X_3345_ _0566_ _1134_ VSS VSS VCC VCC _1135_ sky130_fd_sc_hs__xor2_4
X_3276_ _1070_ _1071_ VSS VSS VCC VCC _1072_ sky130_fd_sc_hs__nand2_2
X_5015_ u_muldiv.dividend\[8\] _2361_ VSS VSS VCC VCC _2369_ sky130_fd_sc_hs__xor2_1
X_5779_ clknet_leaf_21_i_clk _0422_ VSS VSS VCC VCC u_muldiv.outsign sky130_fd_sc_hs__dfxtp_2
X_3130_ _0934_ _0935_ VSS VSS VCC VCC _0936_ sky130_fd_sc_hs__xnor2_4
X_3061_ u_bits.i_op1\[23\] u_bits.i_op1\[22\] _0649_ VSS VSS VCC VCC _0870_
+ sky130_fd_sc_hs__mux2_1
X_3963_ _1635_ VSS VSS VCC VCC _1636_ sky130_fd_sc_hs__buf_2
X_5702_ clknet_leaf_30_i_clk _0345_ VSS VSS VCC VCC u_muldiv.quotient_msk\[16\]
+ sky130_fd_sc_hs__dfxtp_1
X_2914_ _0728_ csr_data\[20\] VSS VSS VCC VCC _0729_ sky130_fd_sc_hs__or2_1
X_3894_ _0791_ i_op1[1] _1596_ VSS VSS VCC VCC _1598_ sky130_fd_sc_hs__mux2_1
X_5633_ clknet_leaf_42_i_clk _0280_ VSS VSS VCC VCC u_muldiv.add_prev\[19\]
+ sky130_fd_sc_hs__dfxtp_1
X_2845_ _0653_ _0654_ _0655_ u_bits.i_op1\[13\] _0658_ _0659_ VSS VSS VCC VCC
+ _0660_ sky130_fd_sc_hs__mux4_1
X_5564_ clknet_leaf_3_i_clk _0211_ VSS VSS VCC VCC u_muldiv.divisor\[45\]
+ sky130_fd_sc_hs__dfxtp_1
X_4515_ _1583_ VSS VSS VCC VCC _1989_ sky130_fd_sc_hs__clkbuf_4
X_2776_ _0460_ u_bits.i_op2\[9\] u_bits.i_op1\[9\] _0464_ VSS VSS VCC VCC
+ _0591_ sky130_fd_sc_hs__a22o_1
X_5495_ clknet_leaf_43_i_clk _0143_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[13\]
+ sky130_fd_sc_hs__dfxtp_1
X_4446_ u_muldiv.divisor\[55\] _1878_ _1829_ u_muldiv.divisor\[56\] _1945_ VSS VSS
+ VCC VCC _0221_ sky130_fd_sc_hs__o221a_1
X_4377_ _1889_ _1890_ VSS VSS VCC VCC _1891_ sky130_fd_sc_hs__nor2_1
X_3328_ _0629_ _1115_ _0955_ VSS VSS VCC VCC _1121_ sky130_fd_sc_hs__a21oi_1
X_3259_ _0697_ u_bits.i_op1\[28\] _0778_ VSS VSS VCC VCC _1056_ sky130_fd_sc_hs__mux2_1
X_5280_ _0620_ _2610_ _2375_ _0702_ VSS VSS VCC VCC _2611_ sky130_fd_sc_hs__o211a_1
X_4300_ _1171_ _1638_ VSS VSS VCC VCC _1825_ sky130_fd_sc_hs__nor2_1
X_4231_ _0446_ i_csr_read _1789_ VSS VSS VCC VCC _1790_ sky130_fd_sc_hs__mux2_1
X_4162_ _1753_ VSS VSS VCC VCC _0129_ sky130_fd_sc_hs__clkbuf_1
X_3113_ _0673_ VSS VSS VCC VCC _0920_ sky130_fd_sc_hs__buf_4
X_4093_ u_pc_sel.i_pc_next\[7\] i_pc_next[7] _1712_ VSS VSS VCC VCC _1719_
+ sky130_fd_sc_hs__mux2_1
X_3044_ _0812_ _0815_ _0810_ VSS VSS VCC VCC _0854_ sky130_fd_sc_hs__a21bo_1
X_4995_ _0786_ _2350_ VSS VSS VCC VCC _2351_ sky130_fd_sc_hs__xnor2_1
X_3946_ _1625_ VSS VSS VCC VCC _0041_ sky130_fd_sc_hs__clkbuf_1
X_3877_ _0993_ _1585_ VSS VSS VCC VCC _0010_ sky130_fd_sc_hs__nor2_1
X_5616_ clknet_leaf_44_i_clk _0263_ VSS VSS VCC VCC u_muldiv.add_prev\[2\]
+ sky130_fd_sc_hs__dfxtp_1
X_2828_ _0642_ VSS VSS VCC VCC _0643_ sky130_fd_sc_hs__clkbuf_4
X_5547_ clknet_leaf_11_i_clk _0195_ VSS VSS VCC VCC csr_data\[31\] sky130_fd_sc_hs__dfxtp_1
X_2759_ _0571_ _0572_ _0573_ VSS VSS VCC VCC _0574_ sky130_fd_sc_hs__o21a_1
X_5478_ clknet_leaf_46_i_clk _0126_ VSS VSS VCC VCC u_mux.i_group_mux sky130_fd_sc_hs__dfxtp_2
X_4429_ u_bits.i_op2\[21\] _1931_ VSS VSS VCC VCC _1932_ sky130_fd_sc_hs__xnor2_1
X_4780_ u_muldiv.o_div\[9\] u_muldiv.o_div\[10\] _2186_ VSS VSS VCC VCC _2194_
+ sky130_fd_sc_hs__or3_1
X_3800_ u_muldiv.mul\[47\] _0741_ _1521_ VSS VSS VCC VCC _1522_ sky130_fd_sc_hs__a21oi_1
X_3731_ _1337_ _1339_ _0760_ VSS VSS VCC VCC _1457_ sky130_fd_sc_hs__mux2_1
X_3662_ u_bits.i_op2\[6\] _0786_ _0926_ _1392_ VSS VSS VCC VCC _1393_ sky130_fd_sc_hs__o22a_1
X_3593_ u_muldiv.dividend\[2\] _1326_ _1327_ u_muldiv.o_div\[2\] _0717_ VSS VSS
+ VCC VCC _1328_ sky130_fd_sc_hs__a221o_1
X_5401_ clknet_leaf_51_i_clk _0049_ VSS VSS VCC VCC o_reg_write sky130_fd_sc_hs__dfxtp_2
X_5332_ o_add[1] _1579_ VSS VSS VCC VCC _2627_ sky130_fd_sc_hs__and2_1
X_5263_ _2362_ _2594_ _0699_ VSS VSS VCC VCC _2595_ sky130_fd_sc_hs__a21o_1
X_5194_ _2375_ _2527_ _2529_ _2532_ VSS VSS VCC VCC _2533_ sky130_fd_sc_hs__o31a_1
X_4214_ u_wr_mux.i_reg_data2\[24\] i_reg_data2[24] _1778_ VSS VSS VCC VCC
+ _1781_ sky130_fd_sc_hs__mux2_1
X_4145_ _1744_ VSS VSS VCC VCC _0121_ sky130_fd_sc_hs__clkbuf_1
X_4076_ _1689_ _1708_ _1709_ VSS VSS VCC VCC _0087_ sky130_fd_sc_hs__a21o_1
X_3027_ _0666_ _0676_ _0659_ VSS VSS VCC VCC _0838_ sky130_fd_sc_hs__mux2_1
X_4978_ u_muldiv.dividend\[4\] _2315_ u_muldiv.dividend\[5\] VSS VSS VCC VCC
+ _2335_ sky130_fd_sc_hs__o21ai_1
X_3929_ _1616_ VSS VSS VCC VCC _0033_ sky130_fd_sc_hs__clkbuf_1
X_4901_ u_muldiv.quotient_msk\[11\] _2280_ _2281_ u_muldiv.quotient_msk\[12\] VSS
+ VSS VCC VCC _0340_ sky130_fd_sc_hs__a22o_1
X_4832_ u_muldiv.o_div\[20\] _2235_ _2154_ VSS VSS VCC VCC _2236_ sky130_fd_sc_hs__mux2_1
X_4763_ u_muldiv.o_div\[6\] _2171_ _2180_ _2164_ VSS VSS VCC VCC _0303_ sky130_fd_sc_hs__a22o_1
X_4694_ _2116_ VSS VSS VCC VCC _2117_ sky130_fd_sc_hs__inv_2
X_3714_ _1333_ csr_data\[9\] _1388_ VSS VSS VCC VCC _1442_ sky130_fd_sc_hs__o21ai_1
X_3645_ _1376_ _1257_ _0867_ VSS VSS VCC VCC _1377_ sky130_fd_sc_hs__a21o_1
X_3576_ _1255_ _0794_ _1310_ _1257_ _0651_ _1112_ VSS VSS VCC VCC _1311_ sky130_fd_sc_hs__mux4_1
X_5315_ u_muldiv.divisor\[27\] _1838_ _2617_ u_muldiv.divisor\[28\] VSS VSS VCC
+ VCC _0418_ sky130_fd_sc_hs__a22o_1
X_5246_ u_muldiv.dividend\[28\] _2564_ VSS VSS VCC VCC _2580_ sky130_fd_sc_hs__xor2_1
X_5177_ _2517_ VSS VSS VCC VCC _0380_ sky130_fd_sc_hs__clkbuf_1
X_4128_ o_pc_target[7] i_pc_target[7] _1734_ VSS VSS VCC VCC _1736_ sky130_fd_sc_hs__mux2_1
X_4059_ u_bits.i_op2\[26\] _0905_ _1681_ VSS VSS VCC VCC _1698_ sky130_fd_sc_hs__mux2_1
X_3430_ op_cnt\[1\] op_cnt\[2\] op_cnt\[3\] VSS VSS VCC VCC _1200_ sky130_fd_sc_hs__nand3_1
X_3361_ _0568_ _0576_ _0598_ VSS VSS VCC VCC _1146_ sky130_fd_sc_hs__nand3_1
X_5100_ _2040_ _2436_ VSS VSS VCC VCC _2447_ sky130_fd_sc_hs__nand2_1
X_5031_ _2382_ _2383_ VSS VSS VCC VCC _2384_ sky130_fd_sc_hs__xnor2_1
X_3292_ _0617_ _0638_ _1086_ VSS VSS VCC VCC _1087_ sky130_fd_sc_hs__and3_1
X_4815_ _2170_ u_muldiv.o_div\[17\] _2218_ _2196_ VSS VSS VCC VCC _2222_ sky130_fd_sc_hs__a31o_1
X_5795_ clknet_leaf_37_i_clk _0437_ VSS VSS VCC VCC u_muldiv.mul\[43\] sky130_fd_sc_hs__dfxtp_1
X_4746_ _2153_ VSS VSS VCC VCC _2167_ sky130_fd_sc_hs__clkbuf_4
X_4677_ _2033_ _2099_ VSS VSS VCC VCC _2100_ sky130_fd_sc_hs__nand2_1
X_3628_ _0687_ _1360_ VSS VSS VCC VCC _1361_ sky130_fd_sc_hs__nor2_1
X_3559_ _1112_ _0791_ _1293_ _1294_ VSS VSS VCC VCC _1295_ sky130_fd_sc_hs__a2bb2o_1
X_5229_ u_muldiv.dividend\[27\] u_muldiv.dividend\[26\] _2552_ VSS VSS VCC VCC
+ _2564_ sky130_fd_sc_hs__or3_1
X_2930_ _0722_ VSS VSS VCC VCC _0743_ sky130_fd_sc_hs__buf_2
X_4600_ op_cnt\[4\] _2021_ _2024_ VSS VSS VCC VCC _0296_ sky130_fd_sc_hs__o21a_1
X_2861_ u_bits.i_op1\[4\] u_bits.i_op1\[3\] _0656_ VSS VSS VCC VCC _0676_
+ sky130_fd_sc_hs__mux2_1
X_5580_ clknet_leaf_9_i_clk _0227_ VSS VSS VCC VCC u_muldiv.divisor\[61\]
+ sky130_fd_sc_hs__dfxtp_1
X_2792_ _0602_ _0603_ _0590_ _0605_ _0606_ VSS VSS VCC VCC _0607_ sky130_fd_sc_hs__o221a_1
X_4531_ _1997_ VSS VSS VCC VCC _0254_ sky130_fd_sc_hs__clkbuf_1
X_4462_ u_bits.i_op2\[26\] u_bits.i_op2\[27\] _1942_ _1951_ VSS VSS VCC VCC
+ _1958_ sky130_fd_sc_hs__or4_1
X_3413_ _0855_ _0903_ VSS VSS VCC VCC _1184_ sky130_fd_sc_hs__nand2_1
X_4393_ _1487_ _1899_ _1845_ VSS VSS VCC VCC _1903_ sky130_fd_sc_hs__o21a_1
X_3344_ _0571_ _1133_ VSS VSS VCC VCC _1134_ sky130_fd_sc_hs__nand2_1
X_3275_ _1068_ _1069_ VSS VSS VCC VCC _1071_ sky130_fd_sc_hs__or2_1
X_5014_ _2157_ _2359_ _2367_ _2368_ VSS VSS VCC VCC _0366_ sky130_fd_sc_hs__o31a_1
X_5778_ clknet_leaf_8_i_clk _0421_ VSS VSS VCC VCC u_muldiv.divisor\[30\]
+ sky130_fd_sc_hs__dfxtp_1
X_4729_ _1839_ _2135_ _2138_ _2151_ VSS VSS VCC VCC _2152_ sky130_fd_sc_hs__o31a_4
X_3060_ _0692_ u_bits.i_op2\[23\] _0636_ _0868_ VSS VSS VCC VCC _0869_ sky130_fd_sc_hs__o22a_1
X_5701_ clknet_leaf_29_i_clk _0344_ VSS VSS VCC VCC u_muldiv.quotient_msk\[15\]
+ sky130_fd_sc_hs__dfxtp_1
X_3962_ _1204_ _1634_ VSS VSS VCC VCC _1635_ sky130_fd_sc_hs__nor2_4
X_2913_ csr_read VSS VSS VCC VCC _0728_ sky130_fd_sc_hs__clkinv_4
X_3893_ _1597_ VSS VSS VCC VCC _0016_ sky130_fd_sc_hs__clkbuf_1
X_5632_ clknet_leaf_42_i_clk _0279_ VSS VSS VCC VCC u_muldiv.add_prev\[18\]
+ sky130_fd_sc_hs__dfxtp_1
X_2844_ _0533_ VSS VSS VCC VCC _0659_ sky130_fd_sc_hs__clkbuf_4
X_5563_ clknet_leaf_5_i_clk _0210_ VSS VSS VCC VCC u_muldiv.divisor\[44\]
+ sky130_fd_sc_hs__dfxtp_1
X_4514_ _1988_ VSS VSS VCC VCC _0246_ sky130_fd_sc_hs__clkbuf_1
X_2775_ _0584_ _0589_ VSS VSS VCC VCC _0590_ sky130_fd_sc_hs__nand2_1
X_5494_ clknet_leaf_43_i_clk _0142_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[12\]
+ sky130_fd_sc_hs__dfxtp_1
X_4445_ _0905_ _1943_ _1944_ VSS VSS VCC VCC _1945_ sky130_fd_sc_hs__o21ai_1
X_4376_ _1445_ _1852_ _1888_ _1856_ VSS VSS VCC VCC _1890_ sky130_fd_sc_hs__a31o_1
X_3327_ _0914_ _1109_ _1119_ VSS VSS VCC VCC _1120_ sky130_fd_sc_hs__a21o_1
X_3258_ _0920_ _1053_ _1054_ VSS VSS VCC VCC _1055_ sky130_fd_sc_hs__a21bo_1
X_3189_ _0989_ _0990_ VSS VSS VCC VCC _0991_ sky130_fd_sc_hs__nor2_1
Xclkbuf_leaf_13_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_13_i_clk
+ sky130_fd_sc_hs__clkbuf_16
Xclkbuf_leaf_28_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_28_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4230_ _1711_ VSS VSS VCC VCC _1789_ sky130_fd_sc_hs__clkbuf_4
X_4161_ _1274_ i_alu_ctrl[4] _1745_ VSS VSS VCC VCC _1753_ sky130_fd_sc_hs__mux2_1
X_4092_ _1718_ VSS VSS VCC VCC _0094_ sky130_fd_sc_hs__clkbuf_1
X_3112_ _0667_ _0678_ _0758_ VSS VSS VCC VCC _0919_ sky130_fd_sc_hs__mux2_1
X_3043_ _0851_ _0852_ VSS VSS VCC VCC _0853_ sky130_fd_sc_hs__nor2_1
X_4994_ _1310_ _1257_ _2328_ _2292_ VSS VSS VCC VCC _2350_ sky130_fd_sc_hs__o31a_1
X_3945_ _0943_ i_op1[25] _1621_ VSS VSS VCC VCC _1625_ sky130_fd_sc_hs__mux2_1
X_5615_ clknet_leaf_46_i_clk _0262_ VSS VSS VCC VCC u_muldiv.add_prev\[1\]
+ sky130_fd_sc_hs__dfxtp_1
X_3876_ _1587_ VSS VSS VCC VCC _0009_ sky130_fd_sc_hs__clkbuf_1
X_2827_ u_bits.i_op2\[4\] VSS VSS VCC VCC _0642_ sky130_fd_sc_hs__clkbuf_4
X_5546_ clknet_leaf_11_i_clk _0194_ VSS VSS VCC VCC csr_data\[30\] sky130_fd_sc_hs__dfxtp_1
X_2758_ _0564_ _0565_ VSS VSS VCC VCC _0573_ sky130_fd_sc_hs__nand2_1
X_5477_ clknet_leaf_48_i_clk _0125_ VSS VSS VCC VCC u_muldiv.i_is_div sky130_fd_sc_hs__dfxtp_1
X_2689_ _0448_ u_bits.i_op1\[14\] _0497_ _0503_ VSS VSS VCC VCC _0504_ sky130_fd_sc_hs__a31o_1
X_4428_ u_bits.i_op2\[20\] _1927_ _1845_ VSS VSS VCC VCC _1931_ sky130_fd_sc_hs__o21a_1
X_4359_ _1874_ _1875_ VSS VSS VCC VCC _1876_ sky130_fd_sc_hs__nor2_1
X_3730_ _1455_ _1456_ _1336_ u_pc_sel.i_pc_next\[10\] VSS VSS VCC VCC o_result[10]
+ sky130_fd_sc_hs__a2bb2o_2
X_3661_ u_bits.i_op2\[6\] _0786_ _0867_ VSS VSS VCC VCC _1392_ sky130_fd_sc_hs__a21oi_1
X_3592_ _0722_ VSS VSS VCC VCC _1327_ sky130_fd_sc_hs__buf_2
X_5400_ clknet_leaf_1_i_clk _0048_ VSS VSS VCC VCC o_store sky130_fd_sc_hs__dfxtp_2
X_5331_ _2626_ VSS VSS VCC VCC _0425_ sky130_fd_sc_hs__clkbuf_1
X_5262_ _0996_ _1029_ _0697_ _2568_ VSS VSS VCC VCC _2594_ sky130_fd_sc_hs__or4_1
X_5193_ _2288_ _2531_ _1206_ VSS VSS VCC VCC _2532_ sky130_fd_sc_hs__a21oi_1
X_4213_ _1780_ VSS VSS VCC VCC _0153_ sky130_fd_sc_hs__clkbuf_1
X_4144_ o_pc_target[15] i_pc_target[15] _1734_ VSS VSS VCC VCC _1744_ sky130_fd_sc_hs__mux2_1
X_4075_ u_bits.i_op2\[30\] _1634_ _1596_ i_op2[30] VSS VSS VCC VCC _1709_
+ sky130_fd_sc_hs__a22o_1
X_3026_ _0832_ _0833_ _0835_ _0836_ _0825_ _0707_ VSS VSS VCC VCC _0837_ sky130_fd_sc_hs__mux4_1
X_4977_ _2334_ VSS VSS VCC VCC _0363_ sky130_fd_sc_hs__clkbuf_1
X_3928_ _0647_ i_op1[17] _1610_ VSS VSS VCC VCC _1616_ sky130_fd_sc_hs__mux2_1
X_3859_ _0749_ o_add[19] _1575_ _1576_ _0453_ VSS VSS VCC VCC _1577_ sky130_fd_sc_hs__a221o_1
X_5529_ clknet_leaf_15_i_clk _0177_ VSS VSS VCC VCC csr_data\[13\] sky130_fd_sc_hs__dfxtp_1
X_4900_ u_muldiv.quotient_msk\[10\] _2280_ _2281_ u_muldiv.quotient_msk\[11\] VSS
+ VSS VCC VCC _0339_ sky130_fd_sc_hs__a22o_1
X_4831_ _2208_ _2232_ _2233_ _2234_ VSS VSS VCC VCC _2235_ sky130_fd_sc_hs__a31o_1
X_4762_ _2165_ _2178_ _2179_ _1842_ u_muldiv.quotient_msk\[6\] VSS VSS VCC VCC
+ _2180_ sky130_fd_sc_hs__a32o_1
X_4693_ _2114_ _2115_ VSS VSS VCC VCC _2116_ sky130_fd_sc_hs__or2_1
X_3713_ _0454_ _1437_ _1439_ _1440_ _1357_ VSS VSS VCC VCC _1441_ sky130_fd_sc_hs__o221a_1
X_3644_ u_bits.i_op2\[5\] VSS VSS VCC VCC _1376_ sky130_fd_sc_hs__clkbuf_4
Xclkbuf_2_2__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_2__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3575_ u_bits.i_op1\[4\] VSS VSS VCC VCC _1310_ sky130_fd_sc_hs__buf_4
X_5314_ u_muldiv.divisor\[26\] _1838_ _2617_ u_muldiv.divisor\[27\] VSS VSS VCC
+ VCC _0417_ sky130_fd_sc_hs__a22o_1
X_5245_ _1827_ _2577_ _2578_ _1840_ VSS VSS VCC VCC _2579_ sky130_fd_sc_hs__a31o_1
X_5176_ u_muldiv.dividend\[21\] _2516_ _2485_ VSS VSS VCC VCC _2517_ sky130_fd_sc_hs__mux2_1
X_4127_ _1735_ VSS VSS VCC VCC _0112_ sky130_fd_sc_hs__clkbuf_1
X_4058_ _1689_ _1696_ _1697_ VSS VSS VCC VCC _0081_ sky130_fd_sc_hs__a21o_1
X_3009_ _0533_ _0819_ VSS VSS VCC VCC _0820_ sky130_fd_sc_hs__and2b_1
X_3360_ _1145_ VSS VSS VCC VCC o_add[9] sky130_fd_sc_hs__inv_2
X_5030_ _2051_ _2076_ VSS VSS VCC VCC _2383_ sky130_fd_sc_hs__and2b_1
X_3291_ _0699_ u_bits.i_op2\[30\] VSS VSS VCC VCC _1086_ sky130_fd_sc_hs__nand2_2
X_4814_ _2221_ VSS VSS VCC VCC _0313_ sky130_fd_sc_hs__clkbuf_1
X_5794_ clknet_leaf_35_i_clk _0436_ VSS VSS VCC VCC u_muldiv.mul\[42\] sky130_fd_sc_hs__dfxtp_1
X_4745_ _2165_ u_muldiv.o_div\[3\] _2158_ _1913_ VSS VSS VCC VCC _2166_ sky130_fd_sc_hs__a31o_1
X_4676_ u_muldiv.dividend\[20\] u_muldiv.divisor\[20\] VSS VSS VCC VCC _2099_
+ sky130_fd_sc_hs__or2b_1
X_3627_ _1253_ _1261_ _1259_ _1252_ _0760_ _0879_ VSS VSS VCC VCC _1360_ sky130_fd_sc_hs__mux4_1
X_3558_ _1112_ _0791_ _0866_ VSS VSS VCC VCC _1294_ sky130_fd_sc_hs__a21o_1
X_3489_ o_wdata[2] _1233_ _0799_ u_wr_mux.i_reg_data2\[10\] VSS VSS VCC VCC
+ _1236_ sky130_fd_sc_hs__a22o_1
X_5228_ _2563_ VSS VSS VCC VCC _0385_ sky130_fd_sc_hs__clkbuf_1
X_5159_ _0646_ _2492_ _2385_ VSS VSS VCC VCC _2501_ sky130_fd_sc_hs__o21ai_1
X_2860_ _0650_ _0663_ VSS VSS VCC VCC _0675_ sky130_fd_sc_hs__nor2_1
X_2791_ _0582_ _0583_ VSS VSS VCC VCC _0606_ sky130_fd_sc_hs__nand2_1
X_4530_ u_muldiv.mul\[24\] u_muldiv.mul\[25\] _1989_ VSS VSS VCC VCC _1997_
+ sky130_fd_sc_hs__mux2_1
X_4461_ u_muldiv.divisor\[58\] _1836_ _1946_ u_muldiv.divisor\[59\] _1957_ VSS VSS
+ VCC VCC _0224_ sky130_fd_sc_hs__a221o_1
X_3412_ o_add[20] _1172_ _1173_ _1182_ VSS VSS VCC VCC _1183_ sky130_fd_sc_hs__or4_1
X_4392_ u_muldiv.divisor\[44\] _1867_ _1887_ u_muldiv.divisor\[45\] _1902_ VSS VSS
+ VCC VCC _0210_ sky130_fd_sc_hs__a221o_1
X_3343_ _1131_ _1132_ VSS VSS VCC VCC _1133_ sky130_fd_sc_hs__nand2_2
X_3274_ _1068_ _1069_ VSS VSS VCC VCC _1070_ sky130_fd_sc_hs__nand2_4
X_5013_ u_muldiv.dividend\[7\] _2154_ VSS VSS VCC VCC _2368_ sky130_fd_sc_hs__or2_1
X_5777_ clknet_leaf_11_i_clk _0420_ VSS VSS VCC VCC u_muldiv.divisor\[29\]
+ sky130_fd_sc_hs__dfxtp_1
X_2989_ _0628_ _0767_ _0771_ _0801_ VSS VSS VCC VCC _0802_ sky130_fd_sc_hs__or4_1
X_4728_ _1831_ _2150_ VSS VSS VCC VCC _2151_ sky130_fd_sc_hs__nand2_1
X_4659_ u_muldiv.divisor\[15\] u_muldiv.dividend\[15\] VSS VSS VCC VCC _2082_
+ sky130_fd_sc_hs__or2b_1
X_3961_ _1633_ VSS VSS VCC VCC _1634_ sky130_fd_sc_hs__buf_2
X_5700_ clknet_leaf_29_i_clk _0343_ VSS VSS VCC VCC u_muldiv.quotient_msk\[14\]
+ sky130_fd_sc_hs__dfxtp_1
X_2912_ _0454_ _0716_ _0726_ VSS VSS VCC VCC _0727_ sky130_fd_sc_hs__o21a_1
X_3892_ _0917_ i_op1[0] _1596_ VSS VSS VCC VCC _1597_ sky130_fd_sc_hs__mux2_1
X_2843_ _0657_ VSS VSS VCC VCC _0658_ sky130_fd_sc_hs__buf_4
X_5631_ clknet_leaf_41_i_clk _0278_ VSS VSS VCC VCC u_muldiv.add_prev\[17\]
+ sky130_fd_sc_hs__dfxtp_1
X_2774_ _0587_ _0588_ VSS VSS VCC VCC _0589_ sky130_fd_sc_hs__xor2_4
X_5562_ clknet_leaf_5_i_clk _0209_ VSS VSS VCC VCC u_muldiv.divisor\[43\]
+ sky130_fd_sc_hs__dfxtp_1
X_4513_ u_muldiv.mul\[16\] u_muldiv.mul\[17\] _1978_ VSS VSS VCC VCC _1988_
+ sky130_fd_sc_hs__mux2_1
X_5493_ clknet_leaf_50_i_clk _0141_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[11\]
+ sky130_fd_sc_hs__dfxtp_4
X_4444_ _0905_ _1943_ _1832_ VSS VSS VCC VCC _1944_ sky130_fd_sc_hs__a21oi_1
X_4375_ _1868_ _1888_ _1445_ VSS VSS VCC VCC _1889_ sky130_fd_sc_hs__a21oi_1
X_3326_ _1110_ _1114_ _1118_ _0858_ VSS VSS VCC VCC _1119_ sky130_fd_sc_hs__a211o_1
Xclkbuf_leaf_9_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_9_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3257_ _0760_ _0793_ _0796_ _0673_ VSS VSS VCC VCC _1054_ sky130_fd_sc_hs__a211o_1
X_3188_ _0987_ _0988_ VSS VSS VCC VCC _0990_ sky130_fd_sc_hs__nor2_1
X_4160_ _1752_ VSS VSS VCC VCC _0128_ sky130_fd_sc_hs__clkbuf_1
X_3111_ _0707_ _0917_ VSS VSS VCC VCC _0918_ sky130_fd_sc_hs__nand2_1
X_4091_ u_pc_sel.i_pc_next\[6\] i_pc_next[6] _1712_ VSS VSS VCC VCC _1718_
+ sky130_fd_sc_hs__mux2_1
X_3042_ _0849_ _0850_ VSS VSS VCC VCC _0852_ sky130_fd_sc_hs__nor2_1
X_4993_ _1826_ _2348_ VSS VSS VCC VCC _2349_ sky130_fd_sc_hs__nand2_1
X_3944_ _1624_ VSS VSS VCC VCC _0040_ sky130_fd_sc_hs__clkbuf_1
X_3875_ o_add[26] _1579_ VSS VSS VCC VCC _1587_ sky130_fd_sc_hs__and2_1
X_5614_ clknet_leaf_44_i_clk _0261_ VSS VSS VCC VCC u_muldiv.add_prev\[0\]
+ sky130_fd_sc_hs__dfxtp_1
X_2826_ _0630_ u_bits.i_op2\[20\] _0637_ _0640_ VSS VSS VCC VCC _0641_ sky130_fd_sc_hs__o22ai_1
X_5545_ clknet_leaf_11_i_clk _0193_ VSS VSS VCC VCC csr_data\[29\] sky130_fd_sc_hs__dfxtp_1
X_2757_ _0564_ _0565_ VSS VSS VCC VCC _0572_ sky130_fd_sc_hs__nor2_1
X_5476_ clknet_leaf_23_i_clk _0124_ VSS VSS VCC VCC o_funct3[2] sky130_fd_sc_hs__dfxtp_4
X_2688_ u_mux.i_group_mux u_bits.i_op2\[14\] VSS VSS VCC VCC _0503_ sky130_fd_sc_hs__and2b_1
X_4427_ u_muldiv.divisor\[51\] _1878_ _1833_ _1929_ _1930_ VSS VSS VCC VCC
+ _0217_ sky130_fd_sc_hs__o221a_1
X_4358_ _1406_ _1850_ _1873_ _1856_ VSS VSS VCC VCC _1875_ sky130_fd_sc_hs__a31o_1
X_4289_ _1819_ VSS VSS VCC VCC _0190_ sky130_fd_sc_hs__clkbuf_1
X_3309_ _1101_ _1102_ VSS VSS VCC VCC _1103_ sky130_fd_sc_hs__nand2_1
X_3660_ _1390_ _0826_ _0751_ VSS VSS VCC VCC _1391_ sky130_fd_sc_hs__mux2_1
X_3591_ _0633_ VSS VSS VCC VCC _1326_ sky130_fd_sc_hs__buf_2
X_5330_ o_add[0] _1579_ VSS VSS VCC VCC _2626_ sky130_fd_sc_hs__and2_1
X_5261_ _2593_ VSS VSS VCC VCC _0388_ sky130_fd_sc_hs__clkbuf_1
X_4212_ u_wr_mux.i_reg_data2\[23\] i_reg_data2[23] _1778_ VSS VSS VCC VCC
+ _1780_ sky130_fd_sc_hs__mux2_1
X_5192_ _0692_ _2530_ VSS VSS VCC VCC _2531_ sky130_fd_sc_hs__xnor2_1
X_4143_ _1743_ VSS VSS VCC VCC _0120_ sky130_fd_sc_hs__clkbuf_1
X_4074_ u_bits.i_op2\[31\] u_bits.i_op2\[29\] _1198_ VSS VSS VCC VCC _1708_
+ sky130_fd_sc_hs__mux2_1
X_3025_ _0662_ _0665_ _0779_ VSS VSS VCC VCC _0836_ sky130_fd_sc_hs__mux2_1
Xclkbuf_leaf_12_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_12_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4976_ u_muldiv.dividend\[4\] _2333_ _2244_ VSS VSS VCC VCC _2334_ sky130_fd_sc_hs__mux2_1
X_3927_ _1615_ VSS VSS VCC VCC _0032_ sky130_fd_sc_hs__clkbuf_1
X_3858_ _0908_ _1569_ _0955_ VSS VSS VCC VCC _1576_ sky130_fd_sc_hs__a21oi_1
Xclkbuf_leaf_27_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_27_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3789_ _1510_ _1511_ _0730_ u_pc_sel.i_pc_next\[14\] VSS VSS VCC VCC o_result[14]
+ sky130_fd_sc_hs__a2bb2o_2
X_2809_ _0623_ VSS VSS VCC VCC _0624_ sky130_fd_sc_hs__buf_2
X_5528_ clknet_leaf_13_i_clk _0176_ VSS VSS VCC VCC csr_data\[12\] sky130_fd_sc_hs__dfxtp_1
X_5459_ clknet_leaf_10_i_clk _0107_ VSS VSS VCC VCC o_pc_target[1] sky130_fd_sc_hs__dfxtp_2
X_4830_ u_muldiv.quotient_msk\[20\] u_muldiv.o_div\[20\] _1840_ VSS VSS VCC
+ VCC _2234_ sky130_fd_sc_hs__o21a_1
X_4761_ u_muldiv.o_div\[5\] u_muldiv.o_div\[6\] _2173_ VSS VSS VCC VCC _2179_
+ sky130_fd_sc_hs__or3_1
X_4692_ u_muldiv.dividend\[26\] u_muldiv.divisor\[26\] VSS VSS VCC VCC _2115_
+ sky130_fd_sc_hs__and2b_1
X_3712_ u_muldiv.mul\[9\] _1330_ _1400_ VSS VSS VCC VCC _1440_ sky130_fd_sc_hs__o21ai_1
X_3643_ _1374_ _0766_ _0751_ VSS VSS VCC VCC _1375_ sky130_fd_sc_hs__mux2_1
X_5313_ u_muldiv.divisor\[25\] _2616_ _2617_ u_muldiv.divisor\[26\] VSS VSS VCC
+ VCC _0416_ sky130_fd_sc_hs__a22o_1
X_3574_ _1307_ _1308_ _0779_ VSS VSS VCC VCC _1309_ sky130_fd_sc_hs__mux2_1
X_5244_ _1029_ _2576_ VSS VSS VCC VCC _2578_ sky130_fd_sc_hs__or2_1
X_5175_ _1208_ _2506_ _2507_ _2515_ VSS VSS VCC VCC _2516_ sky130_fd_sc_hs__a31o_1
X_4126_ o_pc_target[6] i_pc_target[6] _1734_ VSS VSS VCC VCC _1735_ sky130_fd_sc_hs__mux2_1
X_4057_ _0905_ _1687_ _1675_ i_op2[24] VSS VSS VCC VCC _1697_ sky130_fd_sc_hs__a22o_1
X_3008_ u_bits.i_op1\[26\] u_bits.i_op1\[27\] _0656_ VSS VSS VCC VCC _0819_
+ sky130_fd_sc_hs__mux2_1
X_4959_ _2059_ _2317_ VSS VSS VCC VCC _2318_ sky130_fd_sc_hs__nand2_1
X_3290_ _0835_ _0836_ _0838_ _0840_ _0669_ _0670_ VSS VSS VCC VCC _1085_ sky130_fd_sc_hs__mux4_1
X_4813_ u_muldiv.o_div\[16\] _2220_ _2154_ VSS VSS VCC VCC _2221_ sky130_fd_sc_hs__mux2_1
X_5793_ clknet_leaf_35_i_clk _0435_ VSS VSS VCC VCC u_muldiv.mul\[41\] sky130_fd_sc_hs__dfxtp_1
X_4744_ _1208_ VSS VSS VCC VCC _2165_ sky130_fd_sc_hs__clkbuf_4
X_4675_ _2039_ _2083_ _2095_ _2097_ VSS VSS VCC VCC _2098_ sky130_fd_sc_hs__o31a_1
X_3626_ _1358_ _1359_ _1336_ u_pc_sel.i_pc_next\[3\] VSS VSS VCC VCC o_result[3]
+ sky130_fd_sc_hs__a2bb2o_2
X_3557_ _0620_ _0635_ VSS VSS VCC VCC _1293_ sky130_fd_sc_hs__or2_1
X_5227_ u_muldiv.dividend\[26\] _2562_ _2485_ VSS VSS VCC VCC _2563_ sky130_fd_sc_hs__mux2_1
X_3488_ _1192_ u_wr_mux.i_reg_data2\[25\] _1235_ VSS VSS VCC VCC o_wdata[25]
+ sky130_fd_sc_hs__a21o_2
X_5158_ _2499_ _2100_ VSS VSS VCC VCC _2500_ sky130_fd_sc_hs__xor2_1
X_5089_ _2043_ _2081_ _2042_ VSS VSS VCC VCC _2437_ sky130_fd_sc_hs__o21a_1
X_4109_ _1727_ VSS VSS VCC VCC _0102_ sky130_fd_sc_hs__clkbuf_1
X_2790_ _0592_ _0593_ _0604_ VSS VSS VCC VCC _0605_ sky130_fd_sc_hs__o21ai_1
X_4460_ u_bits.i_op2\[27\] _1955_ _1956_ VSS VSS VCC VCC _1957_ sky130_fd_sc_hs__o21a_1
X_3411_ o_add[12] o_add[16] _1177_ _1181_ VSS VSS VCC VCC _1182_ sky130_fd_sc_hs__or4b_1
X_4391_ _1900_ _1901_ VSS VSS VCC VCC _1902_ sky130_fd_sc_hs__nor2_1
X_3342_ _0551_ VSS VSS VCC VCC _1132_ sky130_fd_sc_hs__inv_2
X_3273_ u_bits.i_op1\[30\] u_muldiv.add_prev\[30\] _0452_ VSS VSS VCC VCC
+ _1069_ sky130_fd_sc_hs__mux2_1
X_5012_ _1209_ _2360_ _2361_ _2366_ VSS VSS VCC VCC _2367_ sky130_fd_sc_hs__a31o_1
X_5776_ clknet_leaf_11_i_clk _0419_ VSS VSS VCC VCC u_muldiv.divisor\[28\]
+ sky130_fd_sc_hs__dfxtp_1
X_2988_ _0672_ _0790_ _0798_ _0800_ VSS VSS VCC VCC _0801_ sky130_fd_sc_hs__o211a_1
X_4727_ _2146_ _2147_ _2148_ _2149_ VSS VSS VCC VCC _2150_ sky130_fd_sc_hs__or4_1
X_4658_ _2046_ _2047_ _2079_ _2044_ _2080_ VSS VSS VCC VCC _2081_ sky130_fd_sc_hs__o311a_1
X_3609_ _1287_ _0752_ _0659_ VSS VSS VCC VCC _1343_ sky130_fd_sc_hs__mux2_1
X_4589_ _1204_ op_cnt\[0\] VSS VSS VCC VCC _0292_ sky130_fd_sc_hs__nor2_1
X_3960_ i_flush i_reset_n VSS VSS VCC VCC _1633_ sky130_fd_sc_hs__or2b_1
X_2911_ u_muldiv.mul\[20\] _0717_ _0720_ u_muldiv.mul\[52\] _0725_ VSS VSS VCC
+ VCC _0726_ sky130_fd_sc_hs__a221o_1
X_3891_ _1595_ VSS VSS VCC VCC _1596_ sky130_fd_sc_hs__clkbuf_4
X_2842_ _0656_ VSS VSS VCC VCC _0657_ sky130_fd_sc_hs__clkbuf_4
X_5630_ clknet_leaf_41_i_clk _0277_ VSS VSS VCC VCC u_muldiv.add_prev\[16\]
+ sky130_fd_sc_hs__dfxtp_1
X_5561_ clknet_leaf_7_i_clk _0208_ VSS VSS VCC VCC u_muldiv.divisor\[42\]
+ sky130_fd_sc_hs__dfxtp_1
X_2773_ u_bits.i_op1\[10\] u_muldiv.add_prev\[10\] _0449_ VSS VSS VCC VCC
+ _0588_ sky130_fd_sc_hs__mux2_2
X_4512_ _1987_ VSS VSS VCC VCC _0245_ sky130_fd_sc_hs__clkbuf_1
X_5492_ clknet_leaf_50_i_clk _0140_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[10\]
+ sky130_fd_sc_hs__dfxtp_4
X_4443_ _1850_ _1942_ VSS VSS VCC VCC _1943_ sky130_fd_sc_hs__nand2_1
X_4374_ u_bits.i_op2\[9\] _1883_ VSS VSS VCC VCC _1888_ sky130_fd_sc_hs__or2_1
X_3325_ _0711_ _0860_ _0911_ _1117_ VSS VSS VCC VCC _1118_ sky130_fd_sc_hs__a31o_1
X_3256_ _0780_ _0787_ _0758_ VSS VSS VCC VCC _1053_ sky130_fd_sc_hs__mux2_1
X_3187_ _0987_ _0988_ VSS VSS VCC VCC _0989_ sky130_fd_sc_hs__and2_1
X_5759_ clknet_leaf_19_i_clk _0402_ VSS VSS VCC VCC u_muldiv.divisor\[11\]
+ sky130_fd_sc_hs__dfxtp_1
X_3110_ u_bits.i_op1\[0\] VSS VSS VCC VCC _0917_ sky130_fd_sc_hs__buf_4
X_4090_ _1717_ VSS VSS VCC VCC _0093_ sky130_fd_sc_hs__clkbuf_1
X_3041_ _0849_ _0850_ VSS VSS VCC VCC _0851_ sky130_fd_sc_hs__and2_1
X_4992_ _2056_ _2071_ _2072_ VSS VSS VCC VCC _2348_ sky130_fd_sc_hs__or3_1
X_3943_ _0904_ i_op1[24] _1621_ VSS VSS VCC VCC _1624_ sky130_fd_sc_hs__mux2_1
X_3874_ _1586_ VSS VSS VCC VCC _0008_ sky130_fd_sc_hs__clkbuf_1
X_5613_ clknet_leaf_34_i_clk _0260_ VSS VSS VCC VCC u_muldiv.mul\[30\] sky130_fd_sc_hs__dfxtp_1
X_2825_ _0618_ _0639_ _0631_ VSS VSS VCC VCC _0640_ sky130_fd_sc_hs__and3_1
X_5544_ clknet_leaf_16_i_clk _0192_ VSS VSS VCC VCC csr_data\[28\] sky130_fd_sc_hs__dfxtp_1
X_2756_ _0549_ _0550_ VSS VSS VCC VCC _0571_ sky130_fd_sc_hs__nand2_1
X_2687_ _0500_ _0501_ VSS VSS VCC VCC _0502_ sky130_fd_sc_hs__nor2_1
X_5475_ clknet_leaf_6_i_clk _0123_ VSS VSS VCC VCC o_funct3[1] sky130_fd_sc_hs__dfxtp_4
X_4426_ u_muldiv.divisor\[52\] _1829_ VSS VSS VCC VCC _1930_ sky130_fd_sc_hs__or2_1
X_4357_ _1868_ _1873_ _1406_ VSS VSS VCC VCC _1874_ sky130_fd_sc_hs__a21oi_1
X_4288_ csr_data\[26\] i_csr_data[26] _1811_ VSS VSS VCC VCC _1819_ sky130_fd_sc_hs__mux2_1
X_3308_ _1095_ _1100_ VSS VSS VCC VCC _1102_ sky130_fd_sc_hs__or2_1
X_3239_ _1029_ u_bits.i_op2\[28\] _0634_ VSS VSS VCC VCC _1038_ sky130_fd_sc_hs__a21o_1
Xclkbuf_leaf_8_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_8_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3590_ _0719_ VSS VSS VCC VCC _1325_ sky130_fd_sc_hs__buf_2
X_5260_ u_muldiv.dividend\[29\] _2592_ _2485_ VSS VSS VCC VCC _2593_ sky130_fd_sc_hs__mux2_1
X_4211_ _1779_ VSS VSS VCC VCC _0152_ sky130_fd_sc_hs__clkbuf_1
X_5191_ _0768_ _0691_ _2511_ _2292_ VSS VSS VCC VCC _2530_ sky130_fd_sc_hs__o31a_1
X_4142_ o_pc_target[14] i_pc_target[14] _1734_ VSS VSS VCC VCC _1743_ sky130_fd_sc_hs__mux2_1
X_4073_ _1689_ _1706_ _1707_ VSS VSS VCC VCC _0086_ sky130_fd_sc_hs__a21o_1
X_3024_ _0834_ _0661_ _0783_ VSS VSS VCC VCC _0835_ sky130_fd_sc_hs__mux2_1
X_4975_ _2331_ _2332_ _2229_ VSS VSS VCC VCC _2333_ sky130_fd_sc_hs__mux2_1
X_3926_ _0653_ i_op1[16] _1610_ VSS VSS VCC VCC _1615_ sky130_fd_sc_hs__mux2_1
X_3857_ _0858_ _1568_ _1571_ _1574_ VSS VSS VCC VCC _1575_ sky130_fd_sc_hs__or4_1
X_3788_ _1333_ csr_data\[14\] _1388_ VSS VSS VCC VCC _1511_ sky130_fd_sc_hs__o21ai_1
X_2808_ u_mux.i_add_override _0622_ VSS VSS VCC VCC _0623_ sky130_fd_sc_hs__nor2_2
X_5527_ clknet_leaf_13_i_clk _0175_ VSS VSS VCC VCC csr_data\[11\] sky130_fd_sc_hs__dfxtp_1
X_2739_ _0455_ _0553_ VSS VSS VCC VCC _0554_ sky130_fd_sc_hs__xnor2_2
X_5458_ clknet_leaf_50_i_clk _0106_ VSS VSS VCC VCC o_res_src[2] sky130_fd_sc_hs__dfxtp_2
X_5389_ clknet_leaf_49_i_clk _0037_ VSS VSS VCC VCC u_bits.i_op1\[21\] sky130_fd_sc_hs__dfxtp_2
X_4409_ u_bits.i_op2\[17\] _1915_ VSS VSS VCC VCC _1916_ sky130_fd_sc_hs__nand2_1
X_4760_ u_muldiv.o_div\[5\] _2173_ u_muldiv.o_div\[6\] VSS VSS VCC VCC _2178_
+ sky130_fd_sc_hs__o21ai_1
X_4691_ u_muldiv.divisor\[26\] u_muldiv.dividend\[26\] VSS VSS VCC VCC _2114_
+ sky130_fd_sc_hs__and2b_1
X_3711_ u_muldiv.mul\[41\] _1325_ _1438_ VSS VSS VCC VCC _1439_ sky130_fd_sc_hs__a21oi_1
X_3642_ _1282_ _1288_ _1284_ _1281_ _0789_ _0920_ VSS VSS VCC VCC _1374_ sky130_fd_sc_hs__mux4_1
X_5312_ u_muldiv.divisor\[24\] _2616_ _2617_ u_muldiv.divisor\[25\] VSS VSS VCC
+ VCC _0415_ sky130_fd_sc_hs__a22o_1
X_3573_ _0653_ _0647_ _0650_ VSS VSS VCC VCC _1308_ sky130_fd_sc_hs__mux2_1
X_5243_ _1029_ _2576_ VSS VSS VCC VCC _2577_ sky130_fd_sc_hs__nand2_1
X_5174_ _2303_ _2510_ _2514_ VSS VSS VCC VCC _2515_ sky130_fd_sc_hs__a21oi_1
X_4125_ _1711_ VSS VSS VCC VCC _1734_ sky130_fd_sc_hs__clkbuf_4
X_4056_ u_bits.i_op2\[25\] u_bits.i_op2\[23\] _1681_ VSS VSS VCC VCC _1696_
+ sky130_fd_sc_hs__mux2_1
X_3007_ _0691_ _0692_ u_bits.i_op1\[24\] u_bits.i_op1\[25\] _0658_ _0659_ VSS VSS
+ VCC VCC _0818_ sky130_fd_sc_hs__mux4_1
X_4958_ u_muldiv.divisor\[3\] u_muldiv.dividend\[3\] VSS VSS VCC VCC _2317_
+ sky130_fd_sc_hs__or2b_1
X_4889_ u_muldiv.quotient_msk\[1\] _1210_ _2279_ u_muldiv.quotient_msk\[2\] VSS
+ VSS VCC VCC _0330_ sky130_fd_sc_hs__a22o_1
X_3909_ _0785_ i_op1[8] _1599_ VSS VSS VCC VCC _1606_ sky130_fd_sc_hs__mux2_1
Xclkbuf_leaf_11_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_11_i_clk
+ sky130_fd_sc_hs__clkbuf_16
Xclkbuf_leaf_26_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_26_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4812_ _2208_ _2217_ _2218_ _2219_ VSS VSS VCC VCC _2220_ sky130_fd_sc_hs__a31o_1
X_5792_ clknet_leaf_38_i_clk _0434_ VSS VSS VCC VCC u_muldiv.mul\[40\] sky130_fd_sc_hs__dfxtp_1
X_4743_ _2154_ VSS VSS VCC VCC _2164_ sky130_fd_sc_hs__clkbuf_4
X_4674_ _2086_ _2096_ _2094_ VSS VSS VCC VCC _2097_ sky130_fd_sc_hs__or3_1
X_3625_ _1106_ csr_data\[3\] _1124_ VSS VSS VCC VCC _1359_ sky130_fd_sc_hs__o21ai_1
X_3556_ _0920_ _0948_ VSS VSS VCC VCC _1292_ sky130_fd_sc_hs__nand2_1
X_5226_ _2556_ _2561_ _1877_ VSS VSS VCC VCC _2562_ sky130_fd_sc_hs__mux2_1
X_3487_ o_wdata[1] _1233_ _0799_ u_wr_mux.i_reg_data2\[9\] VSS VSS VCC VCC
+ _1235_ sky130_fd_sc_hs__a22o_1
X_5157_ _2036_ _2038_ _2098_ VSS VSS VCC VCC _2499_ sky130_fd_sc_hs__and3_1
X_5088_ _2042_ _2043_ _2081_ VSS VSS VCC VCC _2436_ sky130_fd_sc_hs__or3_1
X_4108_ u_pc_sel.i_pc_next\[14\] i_pc_next[14] _1723_ VSS VSS VCC VCC _1727_
+ sky130_fd_sc_hs__mux2_1
X_4039_ u_bits.i_op2\[20\] u_bits.i_op2\[18\] _1681_ VSS VSS VCC VCC _1684_
+ sky130_fd_sc_hs__mux2_1
X_3410_ _1141_ _1151_ _1180_ VSS VSS VCC VCC _1181_ sky130_fd_sc_hs__and3_1
X_4390_ _1487_ _1852_ _1899_ _1856_ VSS VSS VCC VCC _1901_ sky130_fd_sc_hs__a31o_1
X_3341_ _0528_ _0547_ VSS VSS VCC VCC _1131_ sky130_fd_sc_hs__nor2_1
X_3272_ _0458_ _1067_ VSS VSS VCC VCC _1068_ sky130_fd_sc_hs__xnor2_1
X_5011_ _1880_ _2364_ _2365_ VSS VSS VCC VCC _2366_ sky130_fd_sc_hs__and3_1
X_5775_ clknet_leaf_11_i_clk _0418_ VSS VSS VCC VCC u_muldiv.divisor\[27\]
+ sky130_fd_sc_hs__dfxtp_1
X_2987_ _0625_ _0799_ VSS VSS VCC VCC _0800_ sky130_fd_sc_hs__and2_2
X_4726_ u_muldiv.divisor\[61\] u_muldiv.divisor\[60\] u_muldiv.divisor\[62\] u_muldiv.i_on_end
+ VSS VSS VCC VCC _2149_ sky130_fd_sc_hs__or4_1
X_4657_ u_muldiv.divisor\[13\] u_muldiv.dividend\[13\] VSS VSS VCC VCC _2080_
+ sky130_fd_sc_hs__or2b_1
X_3608_ _1337_ _1339_ _1340_ _1341_ _0789_ _0674_ VSS VSS VCC VCC _1342_ sky130_fd_sc_hs__mux4_1
X_4588_ _2017_ VSS VSS VCC VCC _0291_ sky130_fd_sc_hs__clkbuf_1
X_3539_ _1274_ o_add[0] _0804_ VSS VSS VCC VCC _1276_ sky130_fd_sc_hs__a21oi_1
X_5209_ _2126_ u_muldiv.dividend\[24\] _2540_ _2111_ VSS VSS VCC VCC _2546_
+ sky130_fd_sc_hs__a22o_1
X_2910_ u_muldiv.dividend\[20\] _0721_ _0723_ u_muldiv.o_div\[20\] _0724_ VSS VSS
+ VCC VCC _0725_ sky130_fd_sc_hs__a221o_1
X_3890_ _1594_ VSS VSS VCC VCC _1595_ sky130_fd_sc_hs__buf_4
X_2841_ u_bits.i_op2\[0\] VSS VSS VCC VCC _0656_ sky130_fd_sc_hs__clkbuf_4
X_5560_ clknet_leaf_7_i_clk _0207_ VSS VSS VCC VCC u_muldiv.divisor\[41\]
+ sky130_fd_sc_hs__dfxtp_1
X_2772_ _0456_ _0586_ VSS VSS VCC VCC _0587_ sky130_fd_sc_hs__xnor2_4
X_4511_ u_muldiv.mul\[15\] u_muldiv.mul\[16\] _1978_ VSS VSS VCC VCC _1987_
+ sky130_fd_sc_hs__mux2_1
X_5491_ clknet_leaf_51_i_clk _0139_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[9\]
+ sky130_fd_sc_hs__dfxtp_4
X_4442_ u_bits.i_op2\[22\] u_bits.i_op2\[23\] _1934_ VSS VSS VCC VCC _1942_
+ sky130_fd_sc_hs__or3_1
X_4373_ _1842_ VSS VSS VCC VCC _1887_ sky130_fd_sc_hs__buf_2
X_3324_ _0702_ u_bits.i_op2\[31\] _0636_ _1116_ VSS VSS VCC VCC _1117_ sky130_fd_sc_hs__o22a_1
X_3255_ _0644_ _1051_ _0712_ VSS VSS VCC VCC _1052_ sky130_fd_sc_hs__o21a_1
X_3186_ u_bits.i_op1\[27\] u_muldiv.add_prev\[27\] _0451_ VSS VSS VCC VCC
+ _0988_ sky130_fd_sc_hs__mux2_1
X_5758_ clknet_leaf_19_i_clk _0401_ VSS VSS VCC VCC u_muldiv.divisor\[10\]
+ sky130_fd_sc_hs__dfxtp_1
X_4709_ u_muldiv.divisor\[29\] u_muldiv.dividend\[29\] VSS VSS VCC VCC _2132_
+ sky130_fd_sc_hs__or2b_1
X_5689_ clknet_leaf_26_i_clk _0332_ VSS VSS VCC VCC u_muldiv.quotient_msk\[3\]
+ sky130_fd_sc_hs__dfxtp_1
X_3040_ u_bits.i_op1\[23\] u_muldiv.add_prev\[23\] _0451_ VSS VSS VCC VCC
+ _0850_ sky130_fd_sc_hs__mux2_1
X_4991_ _2056_ _2072_ _2071_ VSS VSS VCC VCC _2347_ sky130_fd_sc_hs__o21a_1
X_3942_ _1623_ VSS VSS VCC VCC _0039_ sky130_fd_sc_hs__clkbuf_1
X_3873_ o_add[25] _1579_ VSS VSS VCC VCC _1586_ sky130_fd_sc_hs__and2_1
X_5612_ clknet_leaf_34_i_clk _0259_ VSS VSS VCC VCC u_muldiv.mul\[29\] sky130_fd_sc_hs__dfxtp_1
X_2824_ _0638_ VSS VSS VCC VCC _0639_ sky130_fd_sc_hs__clkbuf_2
X_5543_ clknet_leaf_16_i_clk _0191_ VSS VSS VCC VCC csr_data\[27\] sky130_fd_sc_hs__dfxtp_1
X_2755_ _0559_ _0560_ VSS VSS VCC VCC _0570_ sky130_fd_sc_hs__nand2_1
X_2686_ u_bits.i_op1\[15\] u_muldiv.add_prev\[15\] _0449_ VSS VSS VCC VCC
+ _0501_ sky130_fd_sc_hs__mux2_1
X_5474_ clknet_leaf_5_i_clk _0122_ VSS VSS VCC VCC o_funct3[0] sky130_fd_sc_hs__dfxtp_4
X_4425_ u_bits.i_op2\[20\] _1928_ VSS VSS VCC VCC _1929_ sky130_fd_sc_hs__xnor2_1
X_4356_ u_bits.i_op2\[4\] _1376_ u_bits.i_op2\[6\] _1859_ VSS VSS VCC VCC
+ _1873_ sky130_fd_sc_hs__or4_1
X_3307_ _1095_ _1100_ VSS VSS VCC VCC _1101_ sky130_fd_sc_hs__nand2_1
X_4287_ _1818_ VSS VSS VCC VCC _0189_ sky130_fd_sc_hs__clkbuf_1
X_3238_ _0858_ _1028_ _1036_ VSS VSS VCC VCC _1037_ sky130_fd_sc_hs__or3_1
X_3169_ _0644_ _0971_ _0712_ VSS VSS VCC VCC _0972_ sky130_fd_sc_hs__o21a_1
X_4210_ u_wr_mux.i_reg_data2\[22\] i_reg_data2[22] _1778_ VSS VSS VCC VCC
+ _1779_ sky130_fd_sc_hs__mux2_1
X_5190_ _2121_ _2528_ VSS VSS VCC VCC _2529_ sky130_fd_sc_hs__and2_1
X_4141_ _1742_ VSS VSS VCC VCC _0119_ sky130_fd_sc_hs__clkbuf_1
X_4072_ u_bits.i_op2\[29\] _1687_ _1596_ i_op2[29] VSS VSS VCC VCC _1707_
+ sky130_fd_sc_hs__a22o_1
X_3023_ _0655_ u_bits.i_op1\[13\] _0658_ VSS VSS VCC VCC _0834_ sky130_fd_sc_hs__mux2_1
X_4974_ u_muldiv.dividend\[4\] _2315_ VSS VSS VCC VCC _2332_ sky130_fd_sc_hs__xor2_1
X_3925_ _1614_ VSS VSS VCC VCC _0031_ sky130_fd_sc_hs__clkbuf_1
X_3856_ _0672_ _1572_ _1573_ _0800_ VSS VSS VCC VCC _1574_ sky130_fd_sc_hs__o211a_1
X_3787_ _1331_ _1506_ _1508_ _1509_ _0728_ VSS VSS VCC VCC _1510_ sky130_fd_sc_hs__o221a_1
X_2807_ _0618_ _0621_ VSS VSS VCC VCC _0622_ sky130_fd_sc_hs__nor2_4
X_5526_ clknet_leaf_15_i_clk _0174_ VSS VSS VCC VCC csr_data\[10\] sky130_fd_sc_hs__dfxtp_1
X_2738_ _0448_ u_bits.i_op1\[7\] _0497_ _0552_ VSS VSS VCC VCC _0553_ sky130_fd_sc_hs__a31o_1
X_5457_ clknet_leaf_8_i_clk _0105_ VSS VSS VCC VCC o_res_src[1] sky130_fd_sc_hs__dfxtp_2
X_2669_ _0480_ _0483_ VSS VSS VCC VCC _0484_ sky130_fd_sc_hs__nand2_1
X_4408_ u_bits.i_op2\[16\] _1910_ _1846_ VSS VSS VCC VCC _1915_ sky130_fd_sc_hs__o21ai_1
X_5388_ clknet_leaf_49_i_clk _0036_ VSS VSS VCC VCC u_bits.i_op1\[20\] sky130_fd_sc_hs__dfxtp_2
X_4339_ u_bits.i_op2\[3\] _0916_ VSS VSS VCC VCC _1859_ sky130_fd_sc_hs__or2_1
X_3710_ u_muldiv.dividend\[9\] _1326_ _1327_ u_muldiv.o_div\[9\] _1383_ VSS VSS
+ VCC VCC _1438_ sky130_fd_sc_hs__a221o_1
X_4690_ u_muldiv.divisor\[27\] u_muldiv.dividend\[27\] VSS VSS VCC VCC _2113_
+ sky130_fd_sc_hs__xnor2_1
X_3641_ _1372_ _1373_ _1336_ u_pc_sel.i_pc_next\[4\] VSS VSS VCC VCC o_result[4]
+ sky130_fd_sc_hs__a2bb2o_2
X_3572_ u_bits.i_op1\[14\] u_bits.i_op1\[15\] _0650_ VSS VSS VCC VCC _1307_
+ sky130_fd_sc_hs__mux2_1
X_5311_ u_muldiv.divisor\[23\] _2616_ _2617_ u_muldiv.divisor\[24\] VSS VSS VCC
+ VCC _0414_ sky130_fd_sc_hs__a22o_1
X_5242_ _0996_ _2568_ _2385_ VSS VSS VCC VCC _2576_ sky130_fd_sc_hs__o21ai_1
X_5173_ _1206_ _2512_ _2513_ _1828_ VSS VSS VCC VCC _2514_ sky130_fd_sc_hs__o31a_1
X_4124_ _1733_ VSS VSS VCC VCC _0111_ sky130_fd_sc_hs__clkbuf_1
X_4055_ _1689_ _1694_ _1695_ VSS VSS VCC VCC _0080_ sky130_fd_sc_hs__a21o_1
X_3006_ u_muldiv.mul\[22\] _0740_ _0741_ u_muldiv.mul\[54\] _0816_ VSS VSS VCC
+ VCC _0817_ sky130_fd_sc_hs__a221o_1
X_4957_ u_muldiv.dividend\[3\] _2301_ VSS VSS VCC VCC _2316_ sky130_fd_sc_hs__nand2_1
X_4888_ _1210_ u_muldiv.quotient_msk\[0\] _2279_ u_muldiv.quotient_msk\[1\] VSS
+ VSS VCC VCC _0329_ sky130_fd_sc_hs__a22o_1
X_3908_ _1605_ VSS VSS VCC VCC _0023_ sky130_fd_sc_hs__clkbuf_1
X_3839_ u_bits.i_op2\[18\] _0645_ _0637_ _1557_ VSS VSS VCC VCC _1558_ sky130_fd_sc_hs__o22a_1
X_5509_ clknet_leaf_50_i_clk _0157_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[27\]
+ sky130_fd_sc_hs__dfxtp_2
Xclkbuf_leaf_7_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_7_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4811_ u_muldiv.quotient_msk\[16\] u_muldiv.o_div\[16\] _1840_ VSS VSS VCC
+ VCC _2219_ sky130_fd_sc_hs__o21a_1
X_5791_ clknet_leaf_38_i_clk _0433_ VSS VSS VCC VCC u_muldiv.mul\[39\] sky130_fd_sc_hs__dfxtp_1
X_4742_ _2157_ _2160_ _2163_ VSS VSS VCC VCC _0299_ sky130_fd_sc_hs__o21a_1
X_4673_ _2087_ _2091_ _2090_ VSS VSS VCC VCC _2096_ sky130_fd_sc_hs__a21o_1
X_3624_ _0454_ _1353_ _1355_ _1356_ _1357_ VSS VSS VCC VCC _1358_ sky130_fd_sc_hs__o221a_1
X_3555_ _1285_ _1290_ _0687_ VSS VSS VCC VCC _1291_ sky130_fd_sc_hs__mux2_1
X_3486_ _1192_ u_wr_mux.i_reg_data2\[24\] _1234_ VSS VSS VCC VCC o_wdata[24]
+ sky130_fd_sc_hs__a21o_2
X_5225_ _2558_ _2560_ _2288_ VSS VSS VCC VCC _2561_ sky130_fd_sc_hs__mux2_1
X_5156_ u_muldiv.dividend\[20\] _2487_ VSS VSS VCC VCC _2498_ sky130_fd_sc_hs__xor2_1
X_5087_ u_muldiv.dividend\[14\] _2423_ VSS VSS VCC VCC _2435_ sky130_fd_sc_hs__xor2_1
X_4107_ _1726_ VSS VSS VCC VCC _0101_ sky130_fd_sc_hs__clkbuf_1
X_4038_ _1665_ _1682_ _1683_ VSS VSS VCC VCC _0075_ sky130_fd_sc_hs__a21o_1
X_3340_ _1130_ VSS VSS VCC VCC o_add[2] sky130_fd_sc_hs__inv_2
X_5010_ _2362_ _2363_ _1258_ VSS VSS VCC VCC _2365_ sky130_fd_sc_hs__a21o_1
X_3271_ _0724_ u_bits.i_op2\[30\] _0465_ u_bits.i_op1\[30\] VSS VSS VCC VCC
+ _1067_ sky130_fd_sc_hs__a22o_1
X_5774_ clknet_leaf_12_i_clk _0417_ VSS VSS VCC VCC u_muldiv.divisor\[26\]
+ sky130_fd_sc_hs__dfxtp_1
X_2986_ _0682_ VSS VSS VCC VCC _0799_ sky130_fd_sc_hs__clkbuf_4
X_4725_ u_muldiv.divisor\[51\] u_muldiv.divisor\[50\] u_muldiv.divisor\[49\] u_muldiv.divisor\[48\]
+ VSS VSS VCC VCC _2148_ sky130_fd_sc_hs__or4_1
X_4656_ _2050_ _2051_ _2077_ _2048_ _2078_ VSS VSS VCC VCC _2079_ sky130_fd_sc_hs__o311a_1
X_3607_ _1258_ _0785_ _1250_ _1305_ _0651_ _0774_ VSS VSS VCC VCC _1341_ sky130_fd_sc_hs__mux4_1
X_4587_ o_add[31] _1584_ VSS VSS VCC VCC _2017_ sky130_fd_sc_hs__and2_1
X_3538_ _1247_ _1264_ _1271_ _1273_ _1274_ VSS VSS VCC VCC _1275_ sky130_fd_sc_hs__a311o_1
X_3469_ _1225_ VSS VSS VCC VCC o_wdata[16] sky130_fd_sc_hs__buf_2
X_5208_ _2545_ VSS VSS VCC VCC _0383_ sky130_fd_sc_hs__clkbuf_1
X_5139_ _2478_ _2480_ _2482_ _2288_ VSS VSS VCC VCC _2483_ sky130_fd_sc_hs__a2bb2o_1
Xclkbuf_leaf_10_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_10_i_clk
+ sky130_fd_sc_hs__clkbuf_16
Xclkbuf_leaf_25_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_25_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_2840_ u_bits.i_op1\[14\] VSS VSS VCC VCC _0655_ sky130_fd_sc_hs__buf_4
X_2771_ _0449_ u_bits.i_op1\[10\] _0497_ _0585_ VSS VSS VCC VCC _0586_ sky130_fd_sc_hs__a31o_1
X_4510_ _1986_ VSS VSS VCC VCC _0244_ sky130_fd_sc_hs__clkbuf_1
X_5490_ clknet_leaf_51_i_clk _0138_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[8\]
+ sky130_fd_sc_hs__dfxtp_4
X_4441_ u_muldiv.divisor\[54\] _1836_ _1887_ u_muldiv.divisor\[55\] _1941_ VSS VSS
+ VCC VCC _0220_ sky130_fd_sc_hs__a221o_1
X_4372_ u_muldiv.divisor\[40\] _1867_ _1843_ u_muldiv.divisor\[41\] _1886_ VSS VSS
+ VCC VCC _0206_ sky130_fd_sc_hs__a221o_1
X_3323_ _0617_ _0638_ _1115_ VSS VSS VCC VCC _1116_ sky130_fd_sc_hs__and3_1
X_3254_ _0670_ _0765_ _0911_ VSS VSS VCC VCC _1051_ sky130_fd_sc_hs__o21a_1
X_3185_ _0458_ _0986_ VSS VSS VCC VCC _0987_ sky130_fd_sc_hs__xnor2_1
X_5757_ clknet_leaf_26_i_clk _0400_ VSS VSS VCC VCC u_muldiv.divisor\[9\]
+ sky130_fd_sc_hs__dfxtp_1
X_2969_ u_bits.i_op1\[15\] u_bits.i_op1\[14\] _0656_ VSS VSS VCC VCC _0782_
+ sky130_fd_sc_hs__mux2_1
X_4708_ _2122_ _2125_ _2129_ _2130_ _2030_ VSS VSS VCC VCC _2131_ sky130_fd_sc_hs__o311ai_4
X_5688_ clknet_leaf_27_i_clk _0331_ VSS VSS VCC VCC u_muldiv.quotient_msk\[2\]
+ sky130_fd_sc_hs__dfxtp_1
X_4639_ u_muldiv.divisor\[1\] u_muldiv.dividend\[1\] VSS VSS VCC VCC _2062_
+ sky130_fd_sc_hs__xnor2_1
X_4990_ u_muldiv.dividend\[6\] _2336_ VSS VSS VCC VCC _2346_ sky130_fd_sc_hs__nand2_1
X_3941_ _0692_ i_op1[23] _1621_ VSS VSS VCC VCC _1623_ sky130_fd_sc_hs__mux2_1
X_3872_ _0903_ _1585_ VSS VSS VCC VCC _0007_ sky130_fd_sc_hs__nor2_1
X_5611_ clknet_leaf_34_i_clk _0258_ VSS VSS VCC VCC u_muldiv.mul\[28\] sky130_fd_sc_hs__dfxtp_1
X_2823_ o_funct3[1] o_funct3[0] VSS VSS VCC VCC _0638_ sky130_fd_sc_hs__nor2_2
X_5542_ clknet_leaf_16_i_clk _0190_ VSS VSS VCC VCC csr_data\[26\] sky130_fd_sc_hs__dfxtp_1
X_2754_ _0554_ _0555_ VSS VSS VCC VCC _0569_ sky130_fd_sc_hs__nor2_1
X_5473_ clknet_leaf_14_i_clk _0121_ VSS VSS VCC VCC o_pc_target[15] sky130_fd_sc_hs__dfxtp_2
X_2685_ _0456_ _0499_ VSS VSS VCC VCC _0500_ sky130_fd_sc_hs__xnor2_1
X_4424_ _1850_ _1927_ VSS VSS VCC VCC _1928_ sky130_fd_sc_hs__nand2_1
X_4355_ u_muldiv.divisor\[37\] _1867_ _1843_ u_muldiv.divisor\[38\] _1872_ VSS VSS
+ VCC VCC _0203_ sky130_fd_sc_hs__a221o_1
X_3306_ _0539_ _1099_ VSS VSS VCC VCC _1100_ sky130_fd_sc_hs__xnor2_1
X_4286_ csr_data\[25\] i_csr_data[25] _1811_ VSS VSS VCC VCC _1818_ sky130_fd_sc_hs__mux2_1
X_3237_ _0925_ _1031_ _1033_ _0914_ _1035_ VSS VSS VCC VCC _1036_ sky130_fd_sc_hs__a221o_1
X_3168_ _0670_ _0970_ _0911_ VSS VSS VCC VCC _0971_ sky130_fd_sc_hs__o21a_1
X_3099_ _0634_ VSS VSS VCC VCC _0906_ sky130_fd_sc_hs__clkbuf_4
X_4140_ o_pc_target[13] i_pc_target[13] _1734_ VSS VSS VCC VCC _1742_ sky130_fd_sc_hs__mux2_1
X_4071_ u_bits.i_op2\[30\] u_bits.i_op2\[28\] _1198_ VSS VSS VCC VCC _1706_
+ sky130_fd_sc_hs__mux2_1
X_3022_ _0645_ _0647_ _0653_ _0654_ _0651_ _0774_ VSS VSS VCC VCC _0833_ sky130_fd_sc_hs__mux4_1
X_4973_ _1826_ _2326_ _2327_ _2329_ _2330_ VSS VSS VCC VCC _2331_ sky130_fd_sc_hs__a32o_1
X_3924_ _0654_ i_op1[15] _1610_ VSS VSS VCC VCC _1614_ sky130_fd_sc_hs__mux2_1
X_3855_ _0687_ _1347_ VSS VSS VCC VCC _1573_ sky130_fd_sc_hs__nand2_1
X_3786_ u_muldiv.mul\[14\] _0748_ _1400_ VSS VSS VCC VCC _1509_ sky130_fd_sc_hs__o21ai_1
X_2806_ _0619_ _0620_ VSS VSS VCC VCC _0621_ sky130_fd_sc_hs__or2_2
X_5525_ clknet_leaf_13_i_clk _0173_ VSS VSS VCC VCC csr_data\[9\] sky130_fd_sc_hs__dfxtp_1
X_2737_ u_mux.i_group_mux u_bits.i_op2\[7\] VSS VSS VCC VCC _0552_ sky130_fd_sc_hs__and2b_1
X_5456_ clknet_leaf_51_i_clk _0104_ VSS VSS VCC VCC o_res_src[0] sky130_fd_sc_hs__dfxtp_2
X_2668_ _0482_ VSS VSS VCC VCC _0483_ sky130_fd_sc_hs__clkinv_2
X_4407_ u_muldiv.divisor\[47\] _1878_ _1829_ u_muldiv.divisor\[48\] _1914_ VSS VSS
+ VCC VCC _0213_ sky130_fd_sc_hs__o221a_1
X_5387_ clknet_leaf_48_i_clk _0035_ VSS VSS VCC VCC u_bits.i_op1\[19\] sky130_fd_sc_hs__dfxtp_2
X_4338_ u_muldiv.divisor\[34\] _1838_ _1843_ u_muldiv.divisor\[35\] _1858_ VSS VSS
+ VCC VCC _0200_ sky130_fd_sc_hs__a221o_1
X_4269_ csr_data\[17\] i_csr_data[17] _1800_ VSS VSS VCC VCC _1809_ sky130_fd_sc_hs__mux2_1
X_3640_ _1106_ csr_data\[4\] _1124_ VSS VSS VCC VCC _1373_ sky130_fd_sc_hs__o21ai_1
X_3571_ _1305_ _1251_ _0777_ _0776_ _0778_ _0783_ VSS VSS VCC VCC _1306_ sky130_fd_sc_hs__mux4_1
X_5310_ u_muldiv.divisor\[22\] _2616_ _2617_ u_muldiv.divisor\[23\] VSS VSS VCC
+ VCC _0413_ sky130_fd_sc_hs__a22o_1
X_5241_ _2303_ _2131_ _2574_ VSS VSS VCC VCC _2575_ sky130_fd_sc_hs__nand3_1
X_5172_ _2295_ _2511_ _0768_ VSS VSS VCC VCC _2513_ sky130_fd_sc_hs__a21oi_1
X_4123_ o_pc_target[5] i_pc_target[5] _1723_ VSS VSS VCC VCC _1733_ sky130_fd_sc_hs__mux2_1
X_4054_ u_bits.i_op2\[23\] _1687_ _1675_ i_op2[23] VSS VSS VCC VCC _1695_
+ sky130_fd_sc_hs__a22o_1
X_3005_ u_muldiv.dividend\[22\] _0742_ _0743_ u_muldiv.o_div\[22\] _0744_ VSS VSS
+ VCC VCC _0816_ sky130_fd_sc_hs__a221o_1
X_4956_ u_muldiv.dividend\[3\] _2301_ VSS VSS VCC VCC _2315_ sky130_fd_sc_hs__or2_1
X_4887_ _1946_ VSS VSS VCC VCC _2279_ sky130_fd_sc_hs__buf_2
X_3907_ _1258_ i_op1[7] _1599_ VSS VSS VCC VCC _1605_ sky130_fd_sc_hs__mux2_1
X_3838_ _0617_ _0639_ _1556_ VSS VSS VCC VCC _1557_ sky130_fd_sc_hs__and3_1
X_5508_ clknet_leaf_50_i_clk _0156_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[26\]
+ sky130_fd_sc_hs__dfxtp_2
X_3769_ _0714_ _1491_ _1492_ _0623_ _1155_ VSS VSS VCC VCC _1493_ sky130_fd_sc_hs__o32a_1
X_5439_ clknet_leaf_0_i_clk _0087_ VSS VSS VCC VCC u_bits.i_op2\[30\] sky130_fd_sc_hs__dfxtp_4
X_4810_ u_muldiv.o_div\[15\] u_muldiv.o_div\[16\] _2210_ VSS VSS VCC VCC _2218_
+ sky130_fd_sc_hs__or3_2
X_5790_ clknet_leaf_38_i_clk _0432_ VSS VSS VCC VCC u_muldiv.mul\[38\] sky130_fd_sc_hs__dfxtp_1
X_4741_ _2161_ _2162_ u_muldiv.o_div\[2\] VSS VSS VCC VCC _2163_ sky130_fd_sc_hs__a21o_1
X_4672_ _2086_ _2093_ _2094_ VSS VSS VCC VCC _2095_ sky130_fd_sc_hs__or3_1
X_3623_ _0728_ VSS VSS VCC VCC _1357_ sky130_fd_sc_hs__buf_2
X_3554_ _0940_ _1289_ _0673_ VSS VSS VCC VCC _1290_ sky130_fd_sc_hs__mux2_1
X_3485_ o_wdata[0] _1233_ _0799_ u_wr_mux.i_reg_data2\[8\] VSS VSS VCC VCC
+ _1234_ sky130_fd_sc_hs__a22o_1
X_5224_ _0689_ _2559_ VSS VSS VCC VCC _2560_ sky130_fd_sc_hs__xnor2_1
X_5155_ _2497_ VSS VSS VCC VCC _0378_ sky130_fd_sc_hs__clkbuf_1
X_5086_ _2434_ VSS VSS VCC VCC _0372_ sky130_fd_sc_hs__clkbuf_1
X_4106_ u_pc_sel.i_pc_next\[13\] i_pc_next[13] _1723_ VSS VSS VCC VCC _1726_
+ sky130_fd_sc_hs__mux2_1
X_4037_ u_bits.i_op2\[18\] _1663_ _1675_ i_op2[18] VSS VSS VCC VCC _1683_
+ sky130_fd_sc_hs__a22o_1
X_4939_ u_muldiv.dividend\[1\] _2299_ _2244_ VSS VSS VCC VCC _2300_ sky130_fd_sc_hs__mux2_1
X_3270_ _0739_ csr_data\[29\] _1066_ _0732_ VSS VSS VCC VCC o_result[29] sky130_fd_sc_hs__o211a_2
X_5773_ clknet_leaf_12_i_clk _0416_ VSS VSS VCC VCC u_muldiv.divisor\[25\]
+ sky130_fd_sc_hs__dfxtp_1
X_4724_ u_muldiv.divisor\[59\] u_muldiv.divisor\[58\] u_muldiv.divisor\[57\] u_muldiv.divisor\[56\]
+ VSS VSS VCC VCC _2147_ sky130_fd_sc_hs__or4_1
X_2985_ _0672_ _0797_ VSS VSS VCC VCC _0798_ sky130_fd_sc_hs__nand2_1
X_4655_ u_muldiv.divisor\[11\] u_muldiv.dividend\[11\] VSS VSS VCC VCC _2078_
+ sky130_fd_sc_hs__or2b_1
Xclkbuf_leaf_6_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_6_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3606_ _0794_ _1310_ _1257_ _0786_ _0651_ _0774_ VSS VSS VCC VCC _1340_ sky130_fd_sc_hs__mux4_1
X_4586_ _2016_ VSS VSS VCC VCC _0290_ sky130_fd_sc_hs__clkbuf_1
X_3537_ u_mux.i_add_override VSS VSS VCC VCC _1274_ sky130_fd_sc_hs__buf_2
X_3468_ o_wdata[0] u_wr_mux.i_reg_data2\[16\] _1224_ VSS VSS VCC VCC _1225_
+ sky130_fd_sc_hs__mux2_1
X_5207_ u_muldiv.dividend\[24\] _2544_ _2485_ VSS VSS VCC VCC _2545_ sky130_fd_sc_hs__mux2_1
X_3399_ _0523_ _0601_ _0608_ VSS VSS VCC VCC _1174_ sky130_fd_sc_hs__nand3_2
X_5138_ _0645_ _2481_ VSS VSS VCC VCC _2482_ sky130_fd_sc_hs__xnor2_1
X_5069_ _0777_ _2417_ _1839_ VSS VSS VCC VCC _2419_ sky130_fd_sc_hs__o21a_1
X_2770_ u_mux.i_group_mux u_bits.i_op2\[10\] VSS VSS VCC VCC _0585_ sky130_fd_sc_hs__and2b_1
X_4440_ _1939_ _1940_ _1833_ VSS VSS VCC VCC _1941_ sky130_fd_sc_hs__a21oi_1
X_4371_ _1884_ _1885_ VSS VSS VCC VCC _1886_ sky130_fd_sc_hs__nor2_1
X_3322_ _0702_ u_bits.i_op2\[31\] VSS VSS VCC VCC _1115_ sky130_fd_sc_hs__nand2_1
X_3253_ u_muldiv.mul\[29\] _0740_ _0720_ u_muldiv.mul\[61\] _1049_ VSS VSS VCC
+ VCC _1050_ sky130_fd_sc_hs__a221o_1
X_3184_ _0461_ u_bits.i_op2\[27\] _0465_ u_bits.i_op1\[27\] VSS VSS VCC VCC
+ _0986_ sky130_fd_sc_hs__a22o_1
X_5756_ clknet_leaf_26_i_clk _0399_ VSS VSS VCC VCC u_muldiv.divisor\[8\]
+ sky130_fd_sc_hs__dfxtp_1
X_2968_ u_bits.i_op1\[17\] u_bits.i_op1\[16\] _0656_ VSS VSS VCC VCC _0781_
+ sky130_fd_sc_hs__mux2_1
X_5687_ clknet_leaf_28_i_clk _0330_ VSS VSS VCC VCC u_muldiv.quotient_msk\[1\]
+ sky130_fd_sc_hs__dfxtp_1
X_4707_ u_muldiv.dividend\[28\] u_muldiv.divisor\[28\] VSS VSS VCC VCC _2130_
+ sky130_fd_sc_hs__or2b_1
X_4638_ _2060_ u_muldiv.dividend\[2\] VSS VSS VCC VCC _2061_ sky130_fd_sc_hs__or2_1
X_2899_ u_mux.i_add_override VSS VSS VCC VCC _0714_ sky130_fd_sc_hs__buf_2
X_4569_ _2010_ VSS VSS VCC VCC _0279_ sky130_fd_sc_hs__clkbuf_1
X_3940_ _1622_ VSS VSS VCC VCC _0038_ sky130_fd_sc_hs__clkbuf_1
X_3871_ _0855_ _1585_ VSS VSS VCC VCC _0006_ sky130_fd_sc_hs__nor2_1
X_5610_ clknet_leaf_33_i_clk _0257_ VSS VSS VCC VCC u_muldiv.mul\[27\] sky130_fd_sc_hs__dfxtp_1
X_2822_ _0636_ VSS VSS VCC VCC _0637_ sky130_fd_sc_hs__buf_2
X_5541_ clknet_leaf_15_i_clk _0189_ VSS VSS VCC VCC csr_data\[25\] sky130_fd_sc_hs__dfxtp_2
X_2753_ _0528_ _0547_ _0567_ VSS VSS VCC VCC _0568_ sky130_fd_sc_hs__or3_2
X_5472_ clknet_leaf_14_i_clk _0120_ VSS VSS VCC VCC o_pc_target[14] sky130_fd_sc_hs__dfxtp_2
X_2684_ _0448_ u_bits.i_op1\[15\] _0497_ _0498_ VSS VSS VCC VCC _0499_ sky130_fd_sc_hs__a31o_1
X_4423_ u_bits.i_op2\[18\] u_bits.i_op2\[19\] _1919_ VSS VSS VCC VCC _1927_
+ sky130_fd_sc_hs__or3_1
X_4354_ _1870_ _1871_ VSS VSS VCC VCC _1872_ sky130_fd_sc_hs__nor2_1
X_3305_ _0452_ u_bits.i_op2\[31\] _1098_ VSS VSS VCC VCC _1099_ sky130_fd_sc_hs__o21ai_1
X_4285_ _1817_ VSS VSS VCC VCC _0188_ sky130_fd_sc_hs__clkbuf_1
X_3236_ _1029_ u_bits.i_op2\[28\] _0636_ _1034_ VSS VSS VCC VCC _1035_ sky130_fd_sc_hs__o22a_1
X_3167_ _0822_ _0823_ _0668_ VSS VSS VCC VCC _0970_ sky130_fd_sc_hs__mux2_1
Xclkbuf_leaf_24_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_24_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3098_ u_bits.i_op2\[24\] VSS VSS VCC VCC _0905_ sky130_fd_sc_hs__clkbuf_4
Xclkbuf_leaf_39_i_clk clknet_2_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_39_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5739_ clknet_leaf_21_i_clk _0382_ VSS VSS VCC VCC u_muldiv.dividend\[23\]
+ sky130_fd_sc_hs__dfxtp_2
X_4070_ _1689_ _1704_ _1705_ VSS VSS VCC VCC _0085_ sky130_fd_sc_hs__a21o_1
X_3021_ _0691_ _0630_ _0768_ _0646_ _0779_ _0831_ VSS VSS VCC VCC _0832_ sky130_fd_sc_hs__mux4_1
X_4972_ _1310_ _2295_ _2328_ _1826_ VSS VSS VCC VCC _2330_ sky130_fd_sc_hs__a31oi_1
X_3923_ _1613_ VSS VSS VCC VCC _0030_ sky130_fd_sc_hs__clkbuf_1
X_3854_ _0872_ _0876_ _0875_ _0880_ _0524_ _0789_ VSS VSS VCC VCC _1572_ sky130_fd_sc_hs__mux4_1
X_2805_ o_funct3[0] VSS VSS VCC VCC _0620_ sky130_fd_sc_hs__buf_4
X_3785_ u_muldiv.mul\[46\] _0741_ _1507_ VSS VSS VCC VCC _1508_ sky130_fd_sc_hs__a21oi_1
X_5524_ clknet_leaf_12_i_clk _0172_ VSS VSS VCC VCC csr_data\[8\] sky130_fd_sc_hs__dfxtp_1
X_2736_ _0549_ _0550_ VSS VSS VCC VCC _0551_ sky130_fd_sc_hs__xnor2_1
X_5455_ clknet_leaf_10_i_clk _0103_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[15\]
+ sky130_fd_sc_hs__dfxtp_1
X_2667_ _0478_ _0481_ VSS VSS VCC VCC _0482_ sky130_fd_sc_hs__nand2_1
X_4406_ _1911_ _1912_ _1913_ VSS VSS VCC VCC _1914_ sky130_fd_sc_hs__o21ai_1
X_5386_ clknet_leaf_48_i_clk _0034_ VSS VSS VCC VCC u_bits.i_op1\[18\] sky130_fd_sc_hs__dfxtp_2
X_4337_ _1855_ _1857_ VSS VSS VCC VCC _1858_ sky130_fd_sc_hs__nor2_1
X_4268_ _1808_ VSS VSS VCC VCC _0180_ sky130_fd_sc_hs__clkbuf_1
X_3219_ _0458_ _1018_ VSS VSS VCC VCC _1019_ sky130_fd_sc_hs__xnor2_1
X_4199_ u_wr_mux.i_reg_data2\[17\] i_reg_data2[17] _1767_ VSS VSS VCC VCC
+ _1773_ sky130_fd_sc_hs__mux2_1
X_3570_ u_bits.i_op1\[10\] VSS VSS VCC VCC _1305_ sky130_fd_sc_hs__clkbuf_4
X_5240_ _2030_ _2130_ _2122_ _2125_ _2129_ VSS VSS VCC VCC _2574_ sky130_fd_sc_hs__a2111o_1
X_5171_ _0768_ _2385_ _2511_ VSS VSS VCC VCC _2512_ sky130_fd_sc_hs__and3_1
X_4122_ _1732_ VSS VSS VCC VCC _0110_ sky130_fd_sc_hs__clkbuf_1
X_4053_ _0905_ u_bits.i_op2\[22\] _1681_ VSS VSS VCC VCC _1694_ sky130_fd_sc_hs__mux2_1
X_3004_ _0812_ _0815_ VSS VSS VCC VCC o_add[22] sky130_fd_sc_hs__xor2_4
X_4955_ _2314_ VSS VSS VCC VCC _0361_ sky130_fd_sc_hs__clkbuf_1
X_3906_ _1604_ VSS VSS VCC VCC _0022_ sky130_fd_sc_hs__clkbuf_1
X_4886_ _2167_ _2276_ _2278_ VSS VSS VCC VCC _0328_ sky130_fd_sc_hs__a21oi_1
X_3837_ u_bits.i_op2\[18\] _0645_ VSS VSS VCC VCC _1556_ sky130_fd_sc_hs__nand2_1
X_3768_ _1487_ _0776_ _0906_ VSS VSS VCC VCC _1492_ sky130_fd_sc_hs__a21oi_2
X_5507_ clknet_leaf_50_i_clk _0155_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[25\]
+ sky130_fd_sc_hs__dfxtp_2
X_2719_ u_mux.i_group_mux _0533_ VSS VSS VCC VCC _0534_ sky130_fd_sc_hs__and2b_1
X_3699_ _0454_ _1424_ _1426_ _1427_ _1357_ VSS VSS VCC VCC _1428_ sky130_fd_sc_hs__o221a_1
X_5438_ clknet_leaf_0_i_clk _0086_ VSS VSS VCC VCC u_bits.i_op2\[29\] sky130_fd_sc_hs__dfxtp_4
X_5369_ clknet_leaf_47_i_clk _0017_ VSS VSS VCC VCC u_bits.i_op1\[1\] sky130_fd_sc_hs__dfxtp_1
X_4740_ _1835_ _2158_ u_muldiv.quotient_msk\[2\] VSS VSS VCC VCC _2162_ sky130_fd_sc_hs__a21o_1
X_4671_ _2037_ _2036_ VSS VSS VCC VCC _2094_ sky130_fd_sc_hs__or2b_1
X_3622_ u_muldiv.mul\[3\] _1330_ _1331_ VSS VSS VCC VCC _1356_ sky130_fd_sc_hs__o21ai_1
X_3553_ _1288_ _0754_ _0696_ VSS VSS VCC VCC _1289_ sky130_fd_sc_hs__mux2_1
X_3484_ _0718_ VSS VSS VCC VCC _1233_ sky130_fd_sc_hs__buf_4
X_5223_ _0943_ _2548_ _2385_ VSS VSS VCC VCC _2559_ sky130_fd_sc_hs__o21ai_1
X_5154_ u_muldiv.dividend\[19\] _2496_ _2485_ VSS VSS VCC VCC _2497_ sky130_fd_sc_hs__mux2_1
X_4105_ _1725_ VSS VSS VCC VCC _0100_ sky130_fd_sc_hs__clkbuf_1
X_5085_ u_muldiv.dividend\[13\] _2433_ _2378_ VSS VSS VCC VCC _2434_ sky130_fd_sc_hs__mux2_1
X_4036_ u_bits.i_op2\[19\] u_bits.i_op2\[17\] _1681_ VSS VSS VCC VCC _1682_
+ sky130_fd_sc_hs__mux2_1
X_4938_ _2208_ _2286_ _2287_ _2298_ VSS VSS VCC VCC _2299_ sky130_fd_sc_hs__a31o_1
X_4869_ u_muldiv.quotient_msk\[28\] u_muldiv.o_div\[28\] _1840_ VSS VSS VCC
+ VCC _2265_ sky130_fd_sc_hs__o21a_1
X_5772_ clknet_leaf_11_i_clk _0415_ VSS VSS VCC VCC u_muldiv.divisor\[24\]
+ sky130_fd_sc_hs__dfxtp_1
X_2984_ _0669_ _0793_ _0796_ _0707_ VSS VSS VCC VCC _0797_ sky130_fd_sc_hs__a211o_1
X_4723_ u_muldiv.divisor\[40\] _2140_ _2145_ VSS VSS VCC VCC _2146_ sky130_fd_sc_hs__or3_1
X_4654_ _2054_ _2055_ _2075_ _2052_ _2076_ VSS VSS VCC VCC _2077_ sky130_fd_sc_hs__o311a_1
X_3605_ _1338_ _1286_ _0779_ VSS VSS VCC VCC _1339_ sky130_fd_sc_hs__mux2_1
X_4585_ o_add[30] _2004_ VSS VSS VCC VCC _2016_ sky130_fd_sc_hs__and2_1
X_3536_ _0831_ _0917_ _1272_ VSS VSS VCC VCC _1273_ sky130_fd_sc_hs__a21oi_1
X_5206_ _2536_ _2543_ _1877_ VSS VSS VCC VCC _2544_ sky130_fd_sc_hs__mux2_1
X_3467_ _0619_ VSS VSS VCC VCC _1224_ sky130_fd_sc_hs__buf_4
X_3398_ o_add[11] o_add[14] o_add[18] VSS VSS VCC VCC _1173_ sky130_fd_sc_hs__or3_1
X_5137_ _0647_ _2469_ _2385_ VSS VSS VCC VCC _2481_ sky130_fd_sc_hs__o21ai_1
X_5068_ _0777_ _2417_ VSS VSS VCC VCC _2418_ sky130_fd_sc_hs__nand2_1
X_4019_ u_bits.i_op2\[14\] u_bits.i_op2\[12\] _1657_ VSS VSS VCC VCC _1670_
+ sky130_fd_sc_hs__mux2_1
X_4370_ u_bits.i_op2\[9\] _1852_ _1883_ _1856_ VSS VSS VCC VCC _1885_ sky130_fd_sc_hs__a31o_1
X_3321_ _0873_ _1113_ _0674_ VSS VSS VCC VCC _1114_ sky130_fd_sc_hs__mux2_1
X_3252_ u_muldiv.dividend\[29\] _0721_ _0723_ u_muldiv.o_div\[29\] _0744_ VSS VSS
+ VCC VCC _1049_ sky130_fd_sc_hs__a221o_1
X_3183_ _0739_ csr_data\[26\] _0985_ _0732_ VSS VSS VCC VCC o_result[26] sky130_fd_sc_hs__o211a_2
X_5755_ clknet_leaf_26_i_clk _0398_ VSS VSS VCC VCC u_muldiv.divisor\[7\]
+ sky130_fd_sc_hs__dfxtp_1
X_2967_ _0776_ _0777_ u_bits.i_op1\[11\] u_bits.i_op1\[10\] _0778_ _0779_ VSS VSS
+ VCC VCC _0780_ sky130_fd_sc_hs__mux4_2
X_5686_ clknet_leaf_28_i_clk _0329_ VSS VSS VCC VCC u_muldiv.quotient_msk\[0\]
+ sky130_fd_sc_hs__dfxtp_1
X_4706_ _2118_ _2128_ VSS VSS VCC VCC _2129_ sky130_fd_sc_hs__nor2_1
X_2898_ _0688_ _0709_ _0712_ VSS VSS VCC VCC _0713_ sky130_fd_sc_hs__o21ai_1
X_4637_ u_muldiv.divisor\[2\] VSS VSS VCC VCC _2060_ sky130_fd_sc_hs__inv_2
X_4568_ o_add[19] _2004_ VSS VSS VCC VCC _2010_ sky130_fd_sc_hs__and2_1
X_4499_ u_muldiv.mul\[9\] u_muldiv.mul\[10\] _1978_ VSS VSS VCC VCC _1981_
+ sky130_fd_sc_hs__mux2_1
X_3519_ _0917_ _0791_ _1255_ _0794_ _0831_ _1112_ VSS VSS VCC VCC _1256_ sky130_fd_sc_hs__mux4_1
Xclkbuf_leaf_5_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_5_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3870_ _1584_ VSS VSS VCC VCC _1585_ sky130_fd_sc_hs__clkbuf_4
X_2821_ _0620_ _0635_ VSS VSS VCC VCC _0636_ sky130_fd_sc_hs__nor2_4
X_5540_ clknet_leaf_15_i_clk _0188_ VSS VSS VCC VCC csr_data\[24\] sky130_fd_sc_hs__dfxtp_1
X_2752_ _0551_ _0562_ _0566_ VSS VSS VCC VCC _0567_ sky130_fd_sc_hs__or3_1
X_5471_ clknet_leaf_14_i_clk _0119_ VSS VSS VCC VCC o_pc_target[13] sky130_fd_sc_hs__dfxtp_2
X_2683_ u_mux.i_group_mux u_bits.i_op2\[15\] VSS VSS VCC VCC _0498_ sky130_fd_sc_hs__and2b_1
X_4422_ u_muldiv.divisor\[50\] _1836_ _1887_ u_muldiv.divisor\[51\] _1926_ VSS VSS
+ VCC VCC _0216_ sky130_fd_sc_hs__a221o_1
X_4353_ u_bits.i_op2\[6\] _1850_ _1869_ _1856_ VSS VSS VCC VCC _1871_ sky130_fd_sc_hs__a31o_1
X_4284_ csr_data\[24\] i_csr_data[24] _1811_ VSS VSS VCC VCC _1817_ sky130_fd_sc_hs__mux2_1
X_3304_ _1096_ _1097_ _0452_ VSS VSS VCC VCC _1098_ sky130_fd_sc_hs__o21ai_1
X_3235_ _1029_ u_bits.i_op2\[28\] _0867_ VSS VSS VCC VCC _1034_ sky130_fd_sc_hs__a21oi_1
X_3166_ u_muldiv.mul\[26\] _0740_ _0741_ u_muldiv.mul\[58\] _0968_ VSS VSS VCC
+ VCC _0969_ sky130_fd_sc_hs__a221o_1
X_3097_ u_bits.i_op1\[24\] VSS VSS VCC VCC _0904_ sky130_fd_sc_hs__clkbuf_4
X_3999_ _1406_ _1637_ _1651_ i_op2[7] VSS VSS VCC VCC _1656_ sky130_fd_sc_hs__a22o_1
X_5738_ clknet_leaf_21_i_clk _0381_ VSS VSS VCC VCC u_muldiv.dividend\[22\]
+ sky130_fd_sc_hs__dfxtp_2
X_5669_ clknet_leaf_29_i_clk _0312_ VSS VSS VCC VCC u_muldiv.o_div\[15\] sky130_fd_sc_hs__dfxtp_1
X_3020_ _0778_ VSS VSS VCC VCC _0831_ sky130_fd_sc_hs__buf_4
X_4971_ _2295_ _2328_ _1310_ VSS VSS VCC VCC _2329_ sky130_fd_sc_hs__a21o_1
X_3922_ _0655_ i_op1[14] _1610_ VSS VSS VCC VCC _1613_ sky130_fd_sc_hs__mux2_1
X_3853_ u_bits.i_op2\[19\] _0646_ _0637_ _1570_ VSS VSS VCC VCC _1571_ sky130_fd_sc_hs__o22a_1
X_2804_ o_funct3[1] VSS VSS VCC VCC _0619_ sky130_fd_sc_hs__buf_4
X_3784_ u_muldiv.dividend\[14\] _0742_ _0743_ u_muldiv.o_div\[14\] _1383_ VSS VSS
+ VCC VCC _1507_ sky130_fd_sc_hs__a221o_1
X_5523_ clknet_leaf_12_i_clk _0171_ VSS VSS VCC VCC csr_data\[7\] sky130_fd_sc_hs__dfxtp_1
X_2735_ u_bits.i_op1\[4\] u_muldiv.add_prev\[4\] _0450_ VSS VSS VCC VCC _0550_
+ sky130_fd_sc_hs__mux2_1
X_5454_ clknet_leaf_10_i_clk _0102_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[14\]
+ sky130_fd_sc_hs__dfxtp_1
X_2666_ _0476_ _0477_ VSS VSS VCC VCC _0481_ sky130_fd_sc_hs__or2_1
X_5385_ clknet_leaf_48_i_clk _0033_ VSS VSS VCC VCC u_bits.i_op1\[17\] sky130_fd_sc_hs__dfxtp_2
X_4405_ _1880_ VSS VSS VCC VCC _1913_ sky130_fd_sc_hs__buf_4
X_4336_ _0909_ _0916_ _1852_ _1856_ VSS VSS VCC VCC _1857_ sky130_fd_sc_hs__a31o_1
X_4267_ csr_data\[16\] i_csr_data[16] _1800_ VSS VSS VCC VCC _1808_ sky130_fd_sc_hs__mux2_1
X_4198_ _1772_ VSS VSS VCC VCC _0146_ sky130_fd_sc_hs__clkbuf_1
X_3218_ _0461_ u_bits.i_op2\[28\] _0465_ u_bits.i_op1\[28\] VSS VSS VCC VCC
+ _1018_ sky130_fd_sc_hs__a22o_1
X_3149_ _0628_ _0942_ _0953_ VSS VSS VCC VCC _0954_ sky130_fd_sc_hs__or3_1
Xclkbuf_leaf_23_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_23_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5170_ u_bits.i_op1\[20\] u_bits.i_op1\[19\] _2492_ VSS VSS VCC VCC _2511_
+ sky130_fd_sc_hs__or3_2
X_4121_ o_pc_target[4] i_pc_target[4] _1723_ VSS VSS VCC VCC _1732_ sky130_fd_sc_hs__mux2_1
Xclkbuf_leaf_38_i_clk clknet_2_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_38_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4052_ _1689_ _1692_ _1693_ VSS VSS VCC VCC _0079_ sky130_fd_sc_hs__a21o_1
X_3003_ _0737_ _0736_ _0814_ VSS VSS VCC VCC _0815_ sky130_fd_sc_hs__o21ai_2
X_4954_ u_muldiv.dividend\[2\] _2313_ _2244_ VSS VSS VCC VCC _2314_ sky130_fd_sc_hs__mux2_1
X_3905_ _0786_ i_op1[6] _1599_ VSS VSS VCC VCC _1604_ sky130_fd_sc_hs__mux2_1
X_4885_ _2161_ _2277_ u_muldiv.o_div\[31\] VSS VSS VCC VCC _2278_ sky130_fd_sc_hs__a21oi_1
X_3836_ _0751_ _1316_ _0711_ VSS VSS VCC VCC _1555_ sky130_fd_sc_hs__o21a_1
X_3767_ _0908_ _1490_ VSS VSS VCC VCC _1491_ sky130_fd_sc_hs__nor2_1
X_5506_ clknet_leaf_50_i_clk _0154_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[24\]
+ sky130_fd_sc_hs__dfxtp_2
X_2718_ u_bits.i_op2\[1\] VSS VSS VCC VCC _0533_ sky130_fd_sc_hs__clkbuf_4
X_3698_ u_muldiv.mul\[8\] _1330_ _1400_ VSS VSS VCC VCC _1427_ sky130_fd_sc_hs__o21ai_1
X_2649_ _0463_ VSS VSS VCC VCC _0464_ sky130_fd_sc_hs__buf_2
X_5437_ clknet_leaf_0_i_clk _0085_ VSS VSS VCC VCC u_bits.i_op2\[28\] sky130_fd_sc_hs__dfxtp_4
X_5368_ clknet_leaf_47_i_clk _0016_ VSS VSS VCC VCC u_bits.i_op1\[0\] sky130_fd_sc_hs__dfxtp_2
X_5299_ u_muldiv.divisor\[13\] _2614_ _2615_ u_muldiv.divisor\[14\] VSS VSS VCC
+ VCC _0404_ sky130_fd_sc_hs__a22o_1
X_4319_ _1841_ VSS VSS VCC VCC _1842_ sky130_fd_sc_hs__buf_4
X_4670_ _2089_ _2092_ VSS VSS VCC VCC _2093_ sky130_fd_sc_hs__or2b_1
X_3621_ u_muldiv.mul\[35\] _1325_ _1354_ VSS VSS VCC VCC _1355_ sky130_fd_sc_hs__a21oi_1
X_3552_ _1286_ _1287_ _0648_ VSS VSS VCC VCC _1288_ sky130_fd_sc_hs__mux2_1
X_3483_ _1232_ VSS VSS VCC VCC o_wdata[23] sky130_fd_sc_hs__buf_2
X_5222_ _2116_ _2557_ VSS VSS VCC VCC _2558_ sky130_fd_sc_hs__xnor2_1
X_5153_ _1208_ _2487_ _2488_ _2491_ _2495_ VSS VSS VCC VCC _2496_ sky130_fd_sc_hs__a32o_1
X_4104_ u_pc_sel.i_pc_next\[12\] i_pc_next[12] _1723_ VSS VSS VCC VCC _1725_
+ sky130_fd_sc_hs__mux2_1
X_5084_ _1208_ _2423_ _2424_ _2432_ VSS VSS VCC VCC _2433_ sky130_fd_sc_hs__a31o_1
X_4035_ _1198_ VSS VSS VCC VCC _1681_ sky130_fd_sc_hs__clkbuf_4
X_4937_ _2229_ _2297_ VSS VSS VCC VCC _2298_ sky130_fd_sc_hs__nor2_1
X_4868_ u_muldiv.o_div\[27\] u_muldiv.o_div\[28\] _2258_ VSS VSS VCC VCC _2264_
+ sky130_fd_sc_hs__or3_2
X_3819_ _1106_ csr_data\[16\] _1539_ _1124_ VSS VSS VCC VCC o_result[16] sky130_fd_sc_hs__o211a_2
X_4799_ u_muldiv.o_div\[13\] _2201_ u_muldiv.o_div\[14\] VSS VSS VCC VCC _2209_
+ sky130_fd_sc_hs__o21ai_1
X_5771_ clknet_leaf_12_i_clk _0414_ VSS VSS VCC VCC u_muldiv.divisor\[23\]
+ sky130_fd_sc_hs__dfxtp_1
X_2983_ _0668_ _0795_ VSS VSS VCC VCC _0796_ sky130_fd_sc_hs__nor2_1
X_4722_ _2141_ _2142_ _2143_ _2144_ VSS VSS VCC VCC _2145_ sky130_fd_sc_hs__or4_1
X_4653_ u_muldiv.divisor\[9\] u_muldiv.dividend\[9\] VSS VSS VCC VCC _2076_
+ sky130_fd_sc_hs__or2b_1
X_3604_ u_bits.i_op1\[15\] _0653_ _0650_ VSS VSS VCC VCC _1338_ sky130_fd_sc_hs__mux2_1
X_4584_ _2015_ VSS VSS VCC VCC _0289_ sky130_fd_sc_hs__clkbuf_1
X_3535_ _0634_ VSS VSS VCC VCC _1272_ sky130_fd_sc_hs__buf_2
X_3466_ _1223_ VSS VSS VCC VCC o_wdata[15] sky130_fd_sc_hs__buf_2
X_5205_ _2303_ _2538_ _2539_ _2541_ _2542_ VSS VSS VCC VCC _2543_ sky130_fd_sc_hs__o32ai_1
X_3397_ o_add[21] o_add[22] o_add[15] o_add[19] VSS VSS VCC VCC _1172_ sky130_fd_sc_hs__or4_1
X_5136_ _1826_ _2479_ VSS VSS VCC VCC _2480_ sky130_fd_sc_hs__nand2_1
X_5067_ _1305_ _1251_ _2394_ _2292_ VSS VSS VCC VCC _2417_ sky130_fd_sc_hs__o31a_1
X_4018_ _1665_ _1668_ _1669_ VSS VSS VCC VCC _0069_ sky130_fd_sc_hs__a21o_1
X_3320_ _1111_ _1056_ _1001_ _0944_ _1112_ _0825_ VSS VSS VCC VCC _1113_ sky130_fd_sc_hs__mux4_1
X_3251_ _1047_ _1048_ VSS VSS VCC VCC o_add[29] sky130_fd_sc_hs__xnor2_4
X_3182_ _0969_ _0984_ _0447_ VSS VSS VCC VCC _0985_ sky130_fd_sc_hs__a21o_1
X_5754_ clknet_leaf_26_i_clk _0397_ VSS VSS VCC VCC u_muldiv.divisor\[6\]
+ sky130_fd_sc_hs__dfxtp_1
X_2966_ _0663_ VSS VSS VCC VCC _0779_ sky130_fd_sc_hs__buf_4
X_4705_ _2108_ _2127_ VSS VSS VCC VCC _2128_ sky130_fd_sc_hs__or2_1
X_5685_ clknet_leaf_36_i_clk _0328_ VSS VSS VCC VCC u_muldiv.o_div\[31\] sky130_fd_sc_hs__dfxtp_1
X_2897_ _0711_ VSS VSS VCC VCC _0712_ sky130_fd_sc_hs__buf_2
X_4636_ u_muldiv.dividend\[3\] u_muldiv.divisor\[3\] VSS VSS VCC VCC _2059_
+ sky130_fd_sc_hs__or2b_1
X_4567_ _2009_ _2007_ VSS VSS VCC VCC _0278_ sky130_fd_sc_hs__nor2_1
X_4498_ _1980_ VSS VSS VCC VCC _0238_ sky130_fd_sc_hs__clkbuf_1
X_3518_ u_bits.i_op1\[2\] VSS VSS VCC VCC _1255_ sky130_fd_sc_hs__clkbuf_4
X_3449_ _1194_ _1213_ _1214_ VSS VSS VCC VCC _1215_ sky130_fd_sc_hs__mux2_1
X_5119_ _2464_ VSS VSS VCC VCC _0375_ sky130_fd_sc_hs__clkbuf_1
X_2820_ _0619_ o_funct3[2] VSS VSS VCC VCC _0635_ sky130_fd_sc_hs__nand2_1
X_2751_ _0564_ _0565_ VSS VSS VCC VCC _0566_ sky130_fd_sc_hs__xnor2_4
X_5470_ clknet_leaf_14_i_clk _0118_ VSS VSS VCC VCC o_pc_target[12] sky130_fd_sc_hs__dfxtp_2
X_2682_ _0462_ VSS VSS VCC VCC _0497_ sky130_fd_sc_hs__buf_2
X_4421_ _1924_ _1925_ _1833_ VSS VSS VCC VCC _1926_ sky130_fd_sc_hs__a21oi_1
X_4352_ _1868_ _1869_ u_bits.i_op2\[6\] VSS VSS VCC VCC _1870_ sky130_fd_sc_hs__a21oi_1
X_4283_ _1816_ VSS VSS VCC VCC _0187_ sky130_fd_sc_hs__clkbuf_1
X_3303_ u_bits.i_op1\[31\] _0497_ _0626_ VSS VSS VCC VCC _1097_ sky130_fd_sc_hs__a21oi_1
X_3234_ _1032_ _0680_ _0524_ VSS VSS VCC VCC _1033_ sky130_fd_sc_hs__mux2_1
X_3165_ u_muldiv.dividend\[26\] _0742_ _0743_ u_muldiv.o_div\[26\] _0744_ VSS VSS
+ VCC VCC _0968_ sky130_fd_sc_hs__a221o_1
X_3096_ _0903_ VSS VSS VCC VCC o_add[24] sky130_fd_sc_hs__inv_2
X_3998_ u_bits.i_op2\[8\] u_bits.i_op2\[6\] _1639_ VSS VSS VCC VCC _1655_
+ sky130_fd_sc_hs__mux2_1
X_5737_ clknet_leaf_17_i_clk _0380_ VSS VSS VCC VCC u_muldiv.dividend\[21\]
+ sky130_fd_sc_hs__dfxtp_2
X_2949_ _0663_ _0703_ VSS VSS VCC VCC _0762_ sky130_fd_sc_hs__nand2_1
X_5668_ clknet_leaf_29_i_clk _0311_ VSS VSS VCC VCC u_muldiv.o_div\[14\] sky130_fd_sc_hs__dfxtp_1
X_4619_ _2040_ _2041_ VSS VSS VCC VCC _2042_ sky130_fd_sc_hs__nand2_1
X_5599_ clknet_leaf_35_i_clk _0246_ VSS VSS VCC VCC u_muldiv.mul\[16\] sky130_fd_sc_hs__dfxtp_1
X_4970_ u_bits.i_op1\[2\] u_bits.i_op1\[3\] _2308_ VSS VSS VCC VCC _2328_
+ sky130_fd_sc_hs__or3_4
X_3921_ _1612_ VSS VSS VCC VCC _0029_ sky130_fd_sc_hs__clkbuf_1
X_3852_ _0617_ _0639_ _1569_ VSS VSS VCC VCC _1570_ sky130_fd_sc_hs__and3_1
X_2803_ _0617_ VSS VSS VCC VCC _0618_ sky130_fd_sc_hs__clkbuf_4
X_5522_ clknet_leaf_12_i_clk _0170_ VSS VSS VCC VCC csr_data\[6\] sky130_fd_sc_hs__dfxtp_1
X_3783_ _0714_ _1504_ _1505_ _0623_ _1163_ VSS VSS VCC VCC _1506_ sky130_fd_sc_hs__o32a_1
X_2734_ _0456_ _0548_ VSS VSS VCC VCC _0549_ sky130_fd_sc_hs__xnor2_1
X_5453_ clknet_leaf_10_i_clk _0101_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[13\]
+ sky130_fd_sc_hs__dfxtp_1
X_2665_ _0479_ _0474_ VSS VSS VCC VCC _0480_ sky130_fd_sc_hs__nor2_2
X_5384_ clknet_leaf_48_i_clk _0032_ VSS VSS VCC VCC u_bits.i_op1\[16\] sky130_fd_sc_hs__dfxtp_2
X_4404_ u_bits.i_op2\[16\] _1846_ _1910_ VSS VSS VCC VCC _1912_ sky130_fd_sc_hs__and3_1
X_4335_ _1831_ VSS VSS VCC VCC _1856_ sky130_fd_sc_hs__buf_2
X_4266_ _1807_ VSS VSS VCC VCC _0179_ sky130_fd_sc_hs__clkbuf_1
X_4197_ u_wr_mux.i_reg_data2\[16\] i_reg_data2[16] _1767_ VSS VSS VCC VCC
+ _1772_ sky130_fd_sc_hs__mux2_1
X_3217_ _1015_ _1016_ VSS VSS VCC VCC _1017_ sky130_fd_sc_hs__nand2_1
X_3148_ _0925_ _0946_ _0949_ _0914_ _0952_ VSS VSS VCC VCC _0953_ sky130_fd_sc_hs__a221o_1
X_3079_ _0750_ o_add[23] _0887_ VSS VSS VCC VCC _0888_ sky130_fd_sc_hs__a21o_1
Xclkbuf_leaf_4_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_4_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4120_ _1731_ VSS VSS VCC VCC _0109_ sky130_fd_sc_hs__clkbuf_1
X_4051_ u_bits.i_op2\[22\] _1687_ _1675_ i_op2[22] VSS VSS VCC VCC _1693_
+ sky130_fd_sc_hs__a22o_1
X_3002_ _0734_ _0735_ _0813_ VSS VSS VCC VCC _0814_ sky130_fd_sc_hs__o21ai_1
X_4953_ _2208_ _2301_ _2302_ _2312_ VSS VSS VCC VCC _2313_ sky130_fd_sc_hs__a31o_1
X_3904_ _1603_ VSS VSS VCC VCC _0021_ sky130_fd_sc_hs__clkbuf_1
X_4884_ u_muldiv.quotient_msk\[31\] _1878_ _2271_ VSS VSS VCC VCC _2277_ sky130_fd_sc_hs__a21o_1
X_3835_ u_muldiv.mul\[18\] _0717_ _0720_ u_muldiv.mul\[50\] _1553_ VSS VSS VCC
+ VCC _1554_ sky130_fd_sc_hs__a221o_1
X_3766_ _1110_ _1055_ _1486_ _1248_ _1489_ VSS VSS VCC VCC _1490_ sky130_fd_sc_hs__a221o_1
X_2717_ _0530_ _0531_ VSS VSS VCC VCC _0532_ sky130_fd_sc_hs__xnor2_1
X_5505_ clknet_leaf_47_i_clk _0153_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[23\]
+ sky130_fd_sc_hs__dfxtp_2
X_3697_ u_muldiv.mul\[40\] _1325_ _1425_ VSS VSS VCC VCC _1426_ sky130_fd_sc_hs__a21oi_1
X_5436_ clknet_leaf_1_i_clk _0084_ VSS VSS VCC VCC u_bits.i_op2\[27\] sky130_fd_sc_hs__dfxtp_4
X_2648_ u_mux.i_group_mux _0462_ VSS VSS VCC VCC _0463_ sky130_fd_sc_hs__and2_1
X_5367_ clknet_leaf_23_i_clk _0015_ VSS VSS VCC VCC u_muldiv.mul\[63\] sky130_fd_sc_hs__dfxtp_1
X_5298_ u_muldiv.divisor\[12\] _2614_ _2615_ u_muldiv.divisor\[13\] VSS VSS VCC
+ VCC _0403_ sky130_fd_sc_hs__a22o_1
X_4318_ _1840_ VSS VSS VCC VCC _1841_ sky130_fd_sc_hs__buf_4
X_4249_ _1798_ VSS VSS VCC VCC _0171_ sky130_fd_sc_hs__clkbuf_1
X_3620_ u_muldiv.dividend\[3\] _1326_ _1327_ u_muldiv.o_div\[3\] _0717_ VSS VSS
+ VCC VCC _1354_ sky130_fd_sc_hs__a221o_1
X_3551_ u_bits.i_op1\[19\] _0630_ _0657_ VSS VSS VCC VCC _1287_ sky130_fd_sc_hs__mux2_1
X_3482_ o_wdata[7] u_wr_mux.i_reg_data2\[23\] _1224_ VSS VSS VCC VCC _1232_
+ sky130_fd_sc_hs__mux2_1
X_5221_ _2120_ _2528_ _2112_ _2128_ VSS VSS VCC VCC _2557_ sky130_fd_sc_hs__o31ai_2
X_5152_ _1827_ _2493_ _2494_ _1840_ VSS VSS VCC VCC _2495_ sky130_fd_sc_hs__a31o_1
X_4103_ _1724_ VSS VSS VCC VCC _0099_ sky130_fd_sc_hs__clkbuf_1
X_5083_ _2426_ _2427_ _2431_ VSS VSS VCC VCC _2432_ sky130_fd_sc_hs__o21a_1
X_4034_ _1665_ _1679_ _1680_ VSS VSS VCC VCC _0074_ sky130_fd_sc_hs__a21o_1
X_4936_ _2288_ _2289_ _2290_ _2294_ _2296_ VSS VSS VCC VCC _2297_ sky130_fd_sc_hs__o32a_1
X_4867_ u_muldiv.o_div\[27\] _2258_ u_muldiv.o_div\[28\] VSS VSS VCC VCC _2263_
+ sky130_fd_sc_hs__o21ai_1
X_3818_ _1527_ _1538_ _0446_ VSS VSS VCC VCC _1539_ sky130_fd_sc_hs__a21o_1
X_4798_ _1207_ VSS VSS VCC VCC _2208_ sky130_fd_sc_hs__buf_4
X_3749_ u_bits.i_op2\[12\] _0777_ _1267_ VSS VSS VCC VCC _1474_ sky130_fd_sc_hs__a21oi_1
X_5419_ clknet_leaf_49_i_clk _0067_ VSS VSS VCC VCC u_bits.i_op2\[10\] sky130_fd_sc_hs__dfxtp_1
Xclkbuf_leaf_22_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_22_i_clk
+ sky130_fd_sc_hs__clkbuf_16
Xclkbuf_leaf_37_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_37_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5770_ clknet_leaf_12_i_clk _0413_ VSS VSS VCC VCC u_muldiv.divisor\[22\]
+ sky130_fd_sc_hs__dfxtp_1
X_2982_ u_bits.i_op1\[5\] u_bits.i_op1\[4\] _0794_ u_bits.i_op1\[2\] _0650_ _0648_
+ VSS VSS VCC VCC _0795_ sky130_fd_sc_hs__mux4_2
X_4721_ _1834_ u_muldiv.dividend\[31\] VSS VSS VCC VCC _2144_ sky130_fd_sc_hs__nor2_1
X_4652_ _2056_ _2071_ _2072_ _2074_ VSS VSS VCC VCC _2075_ sky130_fd_sc_hs__o31a_1
X_3603_ _1251_ _0777_ _0776_ _0655_ _0778_ _0779_ VSS VSS VCC VCC _1337_ sky130_fd_sc_hs__mux4_1
X_4583_ o_add[29] _2004_ VSS VSS VCC VCC _2015_ sky130_fd_sc_hs__and2_1
X_3534_ _1265_ _1266_ _1270_ _0906_ VSS VSS VCC VCC _1271_ sky130_fd_sc_hs__o211a_1
X_3465_ u_wr_mux.i_reg_data2\[15\] o_wdata[7] _0718_ VSS VSS VCC VCC _1223_
+ sky130_fd_sc_hs__mux2_1
X_5204_ _2540_ _2111_ _2303_ VSS VSS VCC VCC _2542_ sky130_fd_sc_hs__o21ai_1
X_3396_ u_adder.i_cmp_inverse VSS VSS VCC VCC _1171_ sky130_fd_sc_hs__clkinv_2
X_5135_ _2096_ _2477_ _2086_ VSS VSS VCC VCC _2479_ sky130_fd_sc_hs__a21o_1
X_5066_ _2047_ _2079_ _2046_ VSS VSS VCC VCC _2416_ sky130_fd_sc_hs__o21ai_1
X_4017_ u_bits.i_op2\[12\] _1663_ _1651_ i_op2[12] VSS VSS VCC VCC _1669_
+ sky130_fd_sc_hs__a22o_1
X_4919_ _1209_ VSS VSS VCC VCC _2284_ sky130_fd_sc_hs__clkbuf_4
X_3250_ _1017_ _1023_ _1021_ VSS VSS VCC VCC _1048_ sky130_fd_sc_hs__a21bo_1
X_3181_ _0750_ o_add[26] _0982_ _0983_ _0804_ VSS VSS VCC VCC _0984_ sky130_fd_sc_hs__a221o_1
X_5753_ clknet_leaf_25_i_clk _0396_ VSS VSS VCC VCC u_muldiv.divisor\[5\]
+ sky130_fd_sc_hs__dfxtp_1
X_4704_ _2126_ u_muldiv.dividend\[24\] _2107_ VSS VSS VCC VCC _2127_ sky130_fd_sc_hs__a21oi_1
X_2965_ _0657_ VSS VSS VCC VCC _0778_ sky130_fd_sc_hs__buf_4
X_5684_ clknet_leaf_36_i_clk _0327_ VSS VSS VCC VCC u_muldiv.o_div\[30\] sky130_fd_sc_hs__dfxtp_1
X_2896_ _0642_ _0703_ _0710_ VSS VSS VCC VCC _0711_ sky130_fd_sc_hs__a21oi_4
X_4635_ u_muldiv.dividend\[4\] u_muldiv.divisor\[4\] VSS VSS VCC VCC _2058_
+ sky130_fd_sc_hs__or2b_1
X_4566_ o_add[18] VSS VSS VCC VCC _2009_ sky130_fd_sc_hs__inv_2
X_3517_ _1252_ _1253_ _0760_ VSS VSS VCC VCC _1254_ sky130_fd_sc_hs__mux2_1
X_4497_ u_muldiv.mul\[8\] u_muldiv.mul\[9\] _1978_ VSS VSS VCC VCC _1980_
+ sky130_fd_sc_hs__mux2_1
X_3448_ _1198_ u_muldiv.i_on_wait VSS VSS VCC VCC _1214_ sky130_fd_sc_hs__nor2_8
X_3379_ _0505_ _0506_ VSS VSS VCC VCC _1159_ sky130_fd_sc_hs__or2_1
X_5118_ u_muldiv.dividend\[16\] _2463_ _2378_ VSS VSS VCC VCC _2464_ sky130_fd_sc_hs__mux2_1
X_5049_ _1878_ _2393_ _2400_ VSS VSS VCC VCC _2401_ sky130_fd_sc_hs__o21a_1
X_2750_ u_bits.i_op1\[5\] u_muldiv.add_prev\[5\] _0450_ VSS VSS VCC VCC _0565_
+ sky130_fd_sc_hs__mux2_2
X_2681_ _0474_ _0478_ _0484_ _0494_ _0495_ VSS VSS VCC VCC _0496_ sky130_fd_sc_hs__o221a_1
X_4420_ u_bits.i_op2\[19\] _1923_ VSS VSS VCC VCC _1925_ sky130_fd_sc_hs__or2_1
X_4351_ _0688_ _1376_ _1859_ VSS VSS VCC VCC _1869_ sky130_fd_sc_hs__or3_1
X_4282_ csr_data\[23\] i_csr_data[23] _1811_ VSS VSS VCC VCC _1816_ sky130_fd_sc_hs__mux2_1
X_3302_ u_bits.i_op1\[31\] _0497_ _0626_ VSS VSS VCC VCC _1096_ sky130_fd_sc_hs__and3_1
X_3233_ _0664_ _0667_ _0696_ VSS VSS VCC VCC _1032_ sky130_fd_sc_hs__mux2_1
X_3164_ _0964_ _0967_ VSS VSS VCC VCC o_add[26] sky130_fd_sc_hs__xor2_4
X_3095_ _0901_ _0902_ VSS VSS VCC VCC _0903_ sky130_fd_sc_hs__nand2_1
X_3997_ _1641_ _1653_ _1654_ VSS VSS VCC VCC _0063_ sky130_fd_sc_hs__a21o_1
X_5736_ clknet_leaf_16_i_clk _0379_ VSS VSS VCC VCC u_muldiv.dividend\[20\]
+ sky130_fd_sc_hs__dfxtp_2
X_2948_ _0697_ _0699_ _0656_ VSS VSS VCC VCC _0761_ sky130_fd_sc_hs__mux2_1
X_5667_ clknet_leaf_29_i_clk _0310_ VSS VSS VCC VCC u_muldiv.o_div\[13\] sky130_fd_sc_hs__dfxtp_1
X_4618_ u_muldiv.dividend\[14\] u_muldiv.divisor\[14\] VSS VSS VCC VCC _2041_
+ sky130_fd_sc_hs__or2b_1
X_2879_ _0668_ _0693_ VSS VSS VCC VCC _0694_ sky130_fd_sc_hs__and2b_1
X_5598_ clknet_leaf_35_i_clk _0245_ VSS VSS VCC VCC u_muldiv.mul\[15\] sky130_fd_sc_hs__dfxtp_1
X_4549_ _1128_ _2006_ VSS VSS VCC VCC _0263_ sky130_fd_sc_hs__nor2_1
X_3920_ _0776_ i_op1[13] _1610_ VSS VSS VCC VCC _1612_ sky130_fd_sc_hs__mux2_1
X_3851_ u_bits.i_op2\[19\] _0646_ VSS VSS VCC VCC _1569_ sky130_fd_sc_hs__nand2_1
X_2802_ o_funct3[2] VSS VSS VCC VCC _0617_ sky130_fd_sc_hs__clkbuf_4
X_3782_ u_bits.i_op2\[14\] _0655_ _0906_ VSS VSS VCC VCC _1505_ sky130_fd_sc_hs__a21oi_1
X_5521_ clknet_leaf_12_i_clk _0169_ VSS VSS VCC VCC csr_data\[5\] sky130_fd_sc_hs__dfxtp_1
X_2733_ _0459_ u_bits.i_op2\[4\] u_bits.i_op1\[4\] _0463_ VSS VSS VCC VCC
+ _0548_ sky130_fd_sc_hs__a22o_1
X_5452_ clknet_leaf_10_i_clk _0100_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[12\]
+ sky130_fd_sc_hs__dfxtp_1
X_2664_ _0472_ _0473_ VSS VSS VCC VCC _0479_ sky130_fd_sc_hs__and2_1
X_5383_ clknet_leaf_48_i_clk _0031_ VSS VSS VCC VCC u_bits.i_op1\[15\] sky130_fd_sc_hs__dfxtp_2
X_4403_ _1868_ _1910_ u_bits.i_op2\[16\] VSS VSS VCC VCC _1911_ sky130_fd_sc_hs__a21oi_1
X_4334_ _0916_ _1850_ _0909_ VSS VSS VCC VCC _1855_ sky130_fd_sc_hs__a21oi_1
X_4265_ csr_data\[15\] i_csr_data[15] _1800_ VSS VSS VCC VCC _1807_ sky130_fd_sc_hs__mux2_1
X_4196_ _1771_ VSS VSS VCC VCC _0145_ sky130_fd_sc_hs__clkbuf_1
X_3216_ _0895_ _0896_ _0900_ _0936_ _1013_ VSS VSS VCC VCC _1016_ sky130_fd_sc_hs__a2111o_1
X_3147_ _0943_ u_bits.i_op2\[25\] _0636_ _0951_ VSS VSS VCC VCC _0952_ sky130_fd_sc_hs__o22a_1
X_3078_ _0747_ _0885_ _0886_ _0453_ VSS VSS VCC VCC _0887_ sky130_fd_sc_hs__a31o_1
X_5719_ clknet_leaf_24_i_clk _0362_ VSS VSS VCC VCC u_muldiv.dividend\[3\]
+ sky130_fd_sc_hs__dfxtp_1
X_4050_ u_bits.i_op2\[23\] u_bits.i_op2\[21\] _1681_ VSS VSS VCC VCC _1692_
+ sky130_fd_sc_hs__mux2_1
X_3001_ _0467_ _0468_ _0734_ _0735_ VSS VSS VCC VCC _0813_ sky130_fd_sc_hs__a22o_1
X_4952_ _2303_ _2307_ _2311_ VSS VSS VCC VCC _2312_ sky130_fd_sc_hs__a21oi_1
X_4883_ u_muldiv.o_div\[31\] _2271_ _1913_ VSS VSS VCC VCC _2276_ sky130_fd_sc_hs__a21o_1
X_3903_ _1257_ i_op1[5] _1599_ VSS VSS VCC VCC _1603_ sky130_fd_sc_hs__mux2_1
X_3834_ u_muldiv.dividend\[18\] _0721_ _0723_ u_muldiv.o_div\[18\] _0724_ VSS VSS
+ VCC VCC _1553_ sky130_fd_sc_hs__a221o_1
X_3765_ _1487_ _0776_ _0926_ _1488_ VSS VSS VCC VCC _1489_ sky130_fd_sc_hs__o22a_1
X_3696_ u_muldiv.dividend\[8\] _1326_ _1327_ u_muldiv.o_div\[8\] _1383_ VSS VSS
+ VCC VCC _1425_ sky130_fd_sc_hs__a221o_1
X_2716_ u_bits.i_op1\[2\] u_muldiv.add_prev\[2\] _0450_ VSS VSS VCC VCC _0531_
+ sky130_fd_sc_hs__mux2_1
X_5504_ clknet_leaf_47_i_clk _0152_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[22\]
+ sky130_fd_sc_hs__dfxtp_2
X_2647_ u_bits.i_op2\[0\] u_bits.i_op2\[31\] u_muldiv.i_is_div VSS VSS VCC VCC
+ _0462_ sky130_fd_sc_hs__mux2_1
X_5435_ clknet_leaf_1_i_clk _0083_ VSS VSS VCC VCC u_bits.i_op2\[26\] sky130_fd_sc_hs__dfxtp_4
X_5366_ clknet_leaf_34_i_clk _0014_ VSS VSS VCC VCC u_muldiv.mul\[62\] sky130_fd_sc_hs__dfxtp_1
X_5297_ u_muldiv.divisor\[11\] _2614_ _2615_ u_muldiv.divisor\[12\] VSS VSS VCC
+ VCC _0402_ sky130_fd_sc_hs__a22o_1
X_4317_ _1839_ _1206_ VSS VSS VCC VCC _1840_ sky130_fd_sc_hs__nor2_8
X_4248_ csr_data\[7\] i_csr_data[7] _1789_ VSS VSS VCC VCC _1798_ sky130_fd_sc_hs__mux2_1
X_4179_ _1762_ VSS VSS VCC VCC _0137_ sky130_fd_sc_hs__clkbuf_1
X_3550_ u_bits.i_op1\[17\] _0645_ _0657_ VSS VSS VCC VCC _1286_ sky130_fd_sc_hs__mux2_1
X_5220_ u_muldiv.dividend\[26\] _2552_ VSS VSS VCC VCC _2556_ sky130_fd_sc_hs__xor2_1
X_3481_ _1231_ VSS VSS VCC VCC o_wdata[22] sky130_fd_sc_hs__buf_2
X_5151_ _2295_ _2492_ _0646_ VSS VSS VCC VCC _2494_ sky130_fd_sc_hs__a21o_1
X_5082_ _1827_ _2429_ _2430_ _1840_ VSS VSS VCC VCC _2431_ sky130_fd_sc_hs__a31o_1
X_4102_ u_pc_sel.i_pc_next\[11\] i_pc_next[11] _1723_ VSS VSS VCC VCC _1724_
+ sky130_fd_sc_hs__mux2_1
X_4033_ u_bits.i_op2\[17\] _1663_ _1675_ i_op2[17] VSS VSS VCC VCC _1680_
+ sky130_fd_sc_hs__a22o_1
Xclkbuf_leaf_3_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_3_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4935_ _0917_ _2295_ _0791_ VSS VSS VCC VCC _2296_ sky130_fd_sc_hs__a21oi_1
X_4866_ _2167_ _2260_ _2262_ VSS VSS VCC VCC _0324_ sky130_fd_sc_hs__a21oi_1
X_4797_ _2181_ _2205_ _2207_ VSS VSS VCC VCC _0310_ sky130_fd_sc_hs__a21oi_1
X_3817_ _0749_ o_add[16] _1536_ _1537_ _0453_ VSS VSS VCC VCC _1538_ sky130_fd_sc_hs__a221o_1
X_3748_ _0687_ _1027_ _1471_ _1472_ VSS VSS VCC VCC _1473_ sky130_fd_sc_hs__a22o_1
X_3679_ _0674_ _0925_ _0882_ _1408_ _0858_ VSS VSS VCC VCC _1409_ sky130_fd_sc_hs__a311o_1
X_5418_ clknet_leaf_51_i_clk _0066_ VSS VSS VCC VCC u_bits.i_op2\[9\] sky130_fd_sc_hs__dfxtp_4
X_5349_ o_add[16] _1214_ VSS VSS VCC VCC _2629_ sky130_fd_sc_hs__and2_1
X_2981_ u_bits.i_op1\[3\] VSS VSS VCC VCC _0794_ sky130_fd_sc_hs__clkbuf_4
X_4720_ u_muldiv.divisor\[47\] u_muldiv.divisor\[46\] u_muldiv.divisor\[45\] u_muldiv.divisor\[44\]
+ VSS VSS VCC VCC _2143_ sky130_fd_sc_hs__or4_1
X_4651_ _2073_ _2056_ VSS VSS VCC VCC _2074_ sky130_fd_sc_hs__nor2_1
X_3602_ _1334_ _1335_ _1336_ u_pc_sel.i_pc_next\[2\] VSS VSS VCC VCC o_result[2]
+ sky130_fd_sc_hs__a2bb2o_2
X_4582_ _1024_ _1579_ VSS VSS VCC VCC _0288_ sky130_fd_sc_hs__nor2_1
X_3533_ _0622_ o_add[0] _1269_ VSS VSS VCC VCC _1270_ sky130_fd_sc_hs__a21oi_1
X_3464_ _1222_ VSS VSS VCC VCC o_wdata[14] sky130_fd_sc_hs__buf_2
X_5203_ _2540_ _2111_ VSS VSS VCC VCC _2541_ sky130_fd_sc_hs__and2_1
X_5134_ _2086_ _2096_ _2477_ VSS VSS VCC VCC _2478_ sky130_fd_sc_hs__and3_1
X_3395_ u_adder.i_cmp_inverse _1169_ VSS VSS VCC VCC _1170_ sky130_fd_sc_hs__xnor2_1
X_5065_ _2046_ _2047_ _2079_ VSS VSS VCC VCC _2415_ sky130_fd_sc_hs__or3_1
X_4016_ _1487_ u_bits.i_op2\[11\] _1657_ VSS VSS VCC VCC _1668_ sky130_fd_sc_hs__mux2_1
X_4918_ u_muldiv.quotient_msk\[26\] _2282_ _2283_ u_muldiv.quotient_msk\[27\] VSS
+ VSS VCC VCC _0355_ sky130_fd_sc_hs__a22o_1
X_4849_ u_muldiv.o_div\[23\] _2241_ u_muldiv.o_div\[24\] VSS VSS VCC VCC _2249_
+ sky130_fd_sc_hs__o21ai_1
X_3180_ _0629_ _0978_ _0955_ VSS VSS VCC VCC _0983_ sky130_fd_sc_hs__a21oi_1
X_5752_ clknet_leaf_25_i_clk _0395_ VSS VSS VCC VCC u_muldiv.divisor\[4\]
+ sky130_fd_sc_hs__dfxtp_1
X_2964_ u_bits.i_op1\[12\] VSS VSS VCC VCC _0777_ sky130_fd_sc_hs__buf_4
X_4703_ u_muldiv.divisor\[24\] VSS VSS VCC VCC _2126_ sky130_fd_sc_hs__inv_2
X_5683_ clknet_leaf_32_i_clk _0326_ VSS VSS VCC VCC u_muldiv.o_div\[29\] sky130_fd_sc_hs__dfxtp_1
X_2895_ _0617_ _0682_ VSS VSS VCC VCC _0710_ sky130_fd_sc_hs__nand2_2
X_4634_ u_muldiv.dividend\[5\] u_muldiv.divisor\[5\] VSS VSS VCC VCC _2057_
+ sky130_fd_sc_hs__and2b_1
X_4565_ _1176_ _2007_ VSS VSS VCC VCC _0277_ sky130_fd_sc_hs__nor2_1
X_3516_ u_bits.i_op1\[12\] u_bits.i_op1\[13\] _0655_ u_bits.i_op1\[15\] _0650_ _0648_
+ VSS VSS VCC VCC _1253_ sky130_fd_sc_hs__mux4_1
Xclkbuf_leaf_21_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_21_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4496_ _1979_ VSS VSS VCC VCC _0237_ sky130_fd_sc_hs__clkbuf_1
X_3447_ i_funct3[0] i_funct3[1] VSS VSS VCC VCC _1213_ sky130_fd_sc_hs__nand2_1
X_3378_ _0508_ _0502_ VSS VSS VCC VCC _1158_ sky130_fd_sc_hs__or2_2
X_5117_ _2457_ _2462_ _1877_ VSS VSS VCC VCC _2463_ sky130_fd_sc_hs__mux2_1
X_5048_ _2375_ _2395_ _2396_ _1207_ _2399_ VSS VSS VCC VCC _2400_ sky130_fd_sc_hs__a311o_1
Xclkbuf_leaf_36_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_36_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_2680_ _0472_ _0473_ VSS VSS VCC VCC _0495_ sky130_fd_sc_hs__nand2_1
X_4350_ _1846_ VSS VSS VCC VCC _1868_ sky130_fd_sc_hs__buf_2
X_3301_ _0702_ u_muldiv.add_prev\[31\] _0452_ VSS VSS VCC VCC _1095_ sky130_fd_sc_hs__mux2_1
X_4281_ _1815_ VSS VSS VCC VCC _0186_ sky130_fd_sc_hs__clkbuf_1
X_3232_ _0652_ _0660_ _1030_ _0922_ _0668_ _0673_ VSS VSS VCC VCC _1031_ sky130_fd_sc_hs__mux4_1
X_3163_ _0901_ _0936_ _0966_ VSS VSS VCC VCC _0967_ sky130_fd_sc_hs__o21ai_4
X_3094_ _0895_ _0896_ _0900_ VSS VSS VCC VCC _0902_ sky130_fd_sc_hs__nand3_1
X_3996_ u_bits.i_op2\[6\] _1637_ _1651_ i_op2[6] VSS VSS VCC VCC _1654_ sky130_fd_sc_hs__a22o_1
X_5735_ clknet_leaf_18_i_clk _0378_ VSS VSS VCC VCC u_muldiv.dividend\[19\]
+ sky130_fd_sc_hs__dfxtp_2
X_2947_ _0696_ VSS VSS VCC VCC _0760_ sky130_fd_sc_hs__buf_4
X_5666_ clknet_leaf_29_i_clk _0309_ VSS VSS VCC VCC u_muldiv.o_div\[12\] sky130_fd_sc_hs__dfxtp_1
X_4617_ u_muldiv.divisor\[14\] u_muldiv.dividend\[14\] VSS VSS VCC VCC _2040_
+ sky130_fd_sc_hs__or2b_1
X_2878_ _0630_ _0691_ u_bits.i_op1\[21\] _0692_ _0533_ _0658_ VSS VSS VCC VCC
+ _0693_ sky130_fd_sc_hs__mux4_1
X_5597_ clknet_leaf_35_i_clk _0244_ VSS VSS VCC VCC u_muldiv.mul\[14\] sky130_fd_sc_hs__dfxtp_1
X_4548_ _1130_ _2006_ VSS VSS VCC VCC _0262_ sky130_fd_sc_hs__nor2_1
X_4479_ u_muldiv.quotient_msk\[31\] _1210_ _1913_ VSS VSS VCC VCC _0229_ sky130_fd_sc_hs__a21o_1
X_3850_ _0751_ _1345_ _0711_ VSS VSS VCC VCC _1568_ sky130_fd_sc_hs__o21a_1
X_2801_ _0470_ _0615_ VSS VSS VCC VCC _0616_ sky130_fd_sc_hs__xnor2_4
X_3781_ _0908_ _1503_ VSS VSS VCC VCC _1504_ sky130_fd_sc_hs__nor2_1
X_5520_ clknet_leaf_13_i_clk _0168_ VSS VSS VCC VCC csr_data\[4\] sky130_fd_sc_hs__dfxtp_1
X_2732_ _0532_ _0544_ _0545_ _0546_ VSS VSS VCC VCC _0547_ sky130_fd_sc_hs__o211a_1
X_5451_ clknet_leaf_9_i_clk _0099_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[11\]
+ sky130_fd_sc_hs__dfxtp_1
X_2663_ _0476_ _0477_ VSS VSS VCC VCC _0478_ sky130_fd_sc_hs__nand2_1
X_5382_ clknet_leaf_48_i_clk _0030_ VSS VSS VCC VCC u_bits.i_op1\[14\] sky130_fd_sc_hs__dfxtp_2
X_4402_ u_bits.i_op2\[15\] _1906_ VSS VSS VCC VCC _1910_ sky130_fd_sc_hs__or2_1
X_4333_ u_muldiv.divisor\[33\] _1838_ _1843_ u_muldiv.divisor\[34\] _1854_ VSS VSS
+ VCC VCC _0199_ sky130_fd_sc_hs__a221o_1
X_4264_ _1806_ VSS VSS VCC VCC _0178_ sky130_fd_sc_hs__clkbuf_1
X_3215_ _0962_ _0990_ _1013_ _0966_ _1014_ VSS VSS VCC VCC _1015_ sky130_fd_sc_hs__o221a_1
X_4195_ u_wr_mux.i_reg_data2\[15\] i_reg_data2[15] _1767_ VSS VSS VCC VCC
+ _1771_ sky130_fd_sc_hs__mux2_1
X_3146_ _0617_ _0639_ _0950_ VSS VSS VCC VCC _0951_ sky130_fd_sc_hs__and3_1
X_3077_ _0692_ u_bits.i_op2\[23\] _0634_ VSS VSS VCC VCC _0886_ sky130_fd_sc_hs__a21o_1
X_5718_ clknet_leaf_24_i_clk _0361_ VSS VSS VCC VCC u_muldiv.dividend\[2\]
+ sky130_fd_sc_hs__dfxtp_1
X_3979_ _0923_ _0831_ _1639_ VSS VSS VCC VCC _1642_ sky130_fd_sc_hs__mux2_1
X_5649_ clknet_leaf_10_i_clk _0293_ VSS VSS VCC VCC op_cnt\[1\] sky130_fd_sc_hs__dfxtp_1
X_3000_ _0810_ _0811_ VSS VSS VCC VCC _0812_ sky130_fd_sc_hs__and2_2
X_4951_ _1206_ _2309_ _2310_ _1828_ VSS VSS VCC VCC _2311_ sky130_fd_sc_hs__o31a_1
X_4882_ _2275_ VSS VSS VCC VCC _0327_ sky130_fd_sc_hs__clkbuf_1
X_3902_ _1602_ VSS VSS VCC VCC _0020_ sky130_fd_sc_hs__clkbuf_1
X_3833_ _1106_ csr_data\[17\] _1552_ _1124_ VSS VSS VCC VCC o_result[17] sky130_fd_sc_hs__o211a_2
X_3764_ _1487_ _0776_ _1267_ VSS VSS VCC VCC _1488_ sky130_fd_sc_hs__a21oi_1
X_2715_ _0456_ _0529_ VSS VSS VCC VCC _0530_ sky130_fd_sc_hs__xnor2_1
X_5503_ clknet_leaf_43_i_clk _0151_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[21\]
+ sky130_fd_sc_hs__dfxtp_1
X_3695_ _1274_ _1422_ _1423_ _0624_ _1147_ VSS VSS VCC VCC _1424_ sky130_fd_sc_hs__o32a_1
X_2646_ _0460_ VSS VSS VCC VCC _0461_ sky130_fd_sc_hs__buf_2
X_5434_ clknet_leaf_1_i_clk _0082_ VSS VSS VCC VCC u_bits.i_op2\[25\] sky130_fd_sc_hs__dfxtp_4
X_5365_ clknet_leaf_39_i_clk _0013_ VSS VSS VCC VCC u_muldiv.mul\[61\] sky130_fd_sc_hs__dfxtp_1
X_5296_ u_muldiv.divisor\[10\] _2614_ _2615_ u_muldiv.divisor\[11\] VSS VSS VCC
+ VCC _0401_ sky130_fd_sc_hs__a22o_1
X_4316_ u_muldiv.on_wait VSS VSS VCC VCC _1839_ sky130_fd_sc_hs__clkinv_4
X_4247_ _1797_ VSS VSS VCC VCC _0170_ sky130_fd_sc_hs__clkbuf_1
X_4178_ o_wdata[7] i_reg_data2[7] _1756_ VSS VSS VCC VCC _1762_ sky130_fd_sc_hs__mux2_1
X_3129_ u_bits.i_op1\[25\] u_muldiv.add_prev\[25\] _0452_ VSS VSS VCC VCC
+ _0935_ sky130_fd_sc_hs__mux2_2
X_3480_ o_wdata[6] u_wr_mux.i_reg_data2\[22\] _1224_ VSS VSS VCC VCC _1231_
+ sky130_fd_sc_hs__mux2_1
X_5150_ _0646_ _2362_ _2492_ VSS VSS VCC VCC _2493_ sky130_fd_sc_hs__nand3_1
X_4101_ _1711_ VSS VSS VCC VCC _1723_ sky130_fd_sc_hs__clkbuf_4
X_5081_ _2385_ _2428_ _0776_ VSS VSS VCC VCC _2430_ sky130_fd_sc_hs__a21o_1
X_4032_ u_bits.i_op2\[18\] u_bits.i_op2\[16\] _1657_ VSS VSS VCC VCC _1679_
+ sky130_fd_sc_hs__mux2_1
X_4934_ _2292_ VSS VSS VCC VCC _2295_ sky130_fd_sc_hs__clkbuf_4
X_4865_ _2161_ _2261_ u_muldiv.o_div\[27\] VSS VSS VCC VCC _2262_ sky130_fd_sc_hs__a21oi_1
X_4796_ _2167_ _2206_ u_muldiv.o_div\[13\] VSS VSS VCC VCC _2207_ sky130_fd_sc_hs__a21oi_1
X_3816_ _0629_ _1530_ _0955_ VSS VSS VCC VCC _1537_ sky130_fd_sc_hs__a21oi_1
X_3747_ _0670_ _0695_ _0642_ VSS VSS VCC VCC _1472_ sky130_fd_sc_hs__a21oi_1
X_3678_ _1406_ _1258_ _0926_ _1407_ VSS VSS VCC VCC _1408_ sky130_fd_sc_hs__o22a_1
X_5417_ clknet_leaf_52_i_clk _0065_ VSS VSS VCC VCC u_bits.i_op2\[8\] sky130_fd_sc_hs__dfxtp_4
X_5348_ _1162_ _2628_ VSS VSS VCC VCC _0440_ sky130_fd_sc_hs__nor2_1
X_5279_ _0699_ _2594_ VSS VSS VCC VCC _2610_ sky130_fd_sc_hs__nor2_1
X_2980_ _0783_ _0792_ VSS VSS VCC VCC _0793_ sky130_fd_sc_hs__or2b_1
X_4650_ u_muldiv.divisor\[7\] u_muldiv.dividend\[7\] VSS VSS VCC VCC _2073_
+ sky130_fd_sc_hs__and2b_1
X_3601_ _0730_ VSS VSS VCC VCC _1336_ sky130_fd_sc_hs__clkbuf_2
X_4581_ _0993_ _2007_ VSS VSS VCC VCC _0287_ sky130_fd_sc_hs__nor2_1
X_3532_ _0831_ _0917_ _0926_ _1268_ VSS VSS VCC VCC _1269_ sky130_fd_sc_hs__o22a_1
X_3463_ u_wr_mux.i_reg_data2\[14\] o_wdata[6] _0718_ VSS VSS VCC VCC _1222_
+ sky130_fd_sc_hs__mux2_1
X_5202_ _2120_ _2528_ VSS VSS VCC VCC _2540_ sky130_fd_sc_hs__nor2_1
X_5133_ _2458_ _2093_ VSS VSS VCC VCC _2477_ sky130_fd_sc_hs__or2_1
X_3394_ _1104_ _1105_ _1167_ _1168_ VSS VSS VCC VCC _1169_ sky130_fd_sc_hs__o31a_1
X_5064_ u_muldiv.dividend\[12\] _2403_ VSS VSS VCC VCC _2414_ sky130_fd_sc_hs__xor2_1
X_4015_ _1665_ _1666_ _1667_ VSS VSS VCC VCC _0068_ sky130_fd_sc_hs__a21o_1
X_4917_ u_muldiv.quotient_msk\[25\] _2282_ _2283_ u_muldiv.quotient_msk\[26\] VSS
+ VSS VCC VCC _0354_ sky130_fd_sc_hs__a22o_1
X_4848_ _2181_ _2246_ _2248_ VSS VSS VCC VCC _0320_ sky130_fd_sc_hs__a21oi_1
X_4779_ u_muldiv.o_div\[9\] _2186_ u_muldiv.o_div\[10\] VSS VSS VCC VCC _2193_
+ sky130_fd_sc_hs__o21ai_1
Xclkbuf_leaf_2_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_2_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5751_ clknet_leaf_25_i_clk _0394_ VSS VSS VCC VCC u_muldiv.divisor\[3\]
+ sky130_fd_sc_hs__dfxtp_1
X_2963_ u_bits.i_op1\[13\] VSS VSS VCC VCC _0776_ sky130_fd_sc_hs__clkbuf_4
X_4702_ _2124_ u_muldiv.divisor\[26\] _2123_ u_muldiv.dividend\[27\] VSS VSS VCC
+ VCC _2125_ sky130_fd_sc_hs__a2bb2o_1
X_5682_ clknet_leaf_32_i_clk _0325_ VSS VSS VCC VCC u_muldiv.o_div\[28\] sky130_fd_sc_hs__dfxtp_1
X_2894_ _0708_ VSS VSS VCC VCC _0709_ sky130_fd_sc_hs__inv_2
X_4633_ u_muldiv.divisor\[6\] u_muldiv.dividend\[6\] VSS VSS VCC VCC _2056_
+ sky130_fd_sc_hs__and2b_1
X_4564_ _2008_ VSS VSS VCC VCC _0276_ sky130_fd_sc_hs__clkbuf_1
X_3515_ _0785_ _1250_ u_bits.i_op1\[10\] _1251_ _0778_ _0783_ VSS VSS VCC VCC
+ _1252_ sky130_fd_sc_hs__mux4_1
X_4495_ u_muldiv.mul\[7\] u_muldiv.mul\[8\] _1978_ VSS VSS VCC VCC _1979_
+ sky130_fd_sc_hs__mux2_1
X_3446_ i_flush _1212_ VSS VSS VCC VCC _0002_ sky130_fd_sc_hs__nor2_1
X_3377_ _1157_ VSS VSS VCC VCC o_add[12] sky130_fd_sc_hs__inv_2
X_5116_ _2459_ _2461_ _2288_ VSS VSS VCC VCC _2462_ sky130_fd_sc_hs__mux2_1
X_5047_ u_muldiv.on_wait _2397_ _2398_ VSS VSS VCC VCC _2399_ sky130_fd_sc_hs__and3_1
X_3300_ _1073_ _1075_ _1076_ _1072_ VSS VSS VCC VCC _1094_ sky130_fd_sc_hs__a31o_2
X_4280_ csr_data\[22\] i_csr_data[22] _1811_ VSS VSS VCC VCC _1815_ sky130_fd_sc_hs__mux2_1
X_3231_ _1029_ u_bits.i_op1\[27\] _0689_ _0943_ _0778_ _0779_ VSS VSS VCC VCC
+ _1030_ sky130_fd_sc_hs__mux4_1
X_3162_ _0934_ _0935_ _0965_ VSS VSS VCC VCC _0966_ sky130_fd_sc_hs__o21ai_2
X_3093_ _0895_ _0896_ _0900_ VSS VSS VCC VCC _0901_ sky130_fd_sc_hs__a21o_1
X_5803_ clknet_leaf_34_i_clk _0445_ VSS VSS VCC VCC u_muldiv.mul\[51\] sky130_fd_sc_hs__dfxtp_1
X_3995_ _1406_ _1376_ _1639_ VSS VSS VCC VCC _1653_ sky130_fd_sc_hs__mux2_1
X_5734_ clknet_leaf_18_i_clk _0377_ VSS VSS VCC VCC u_muldiv.dividend\[18\]
+ sky130_fd_sc_hs__dfxtp_2
X_2946_ _0754_ _0757_ _0758_ VSS VSS VCC VCC _0759_ sky130_fd_sc_hs__mux2_1
X_5665_ clknet_leaf_29_i_clk _0308_ VSS VSS VCC VCC u_muldiv.o_div\[11\] sky130_fd_sc_hs__dfxtp_1
X_2877_ u_bits.i_op1\[23\] VSS VSS VCC VCC _0692_ sky130_fd_sc_hs__clkbuf_4
X_4616_ u_muldiv.dividend\[15\] u_muldiv.divisor\[15\] VSS VSS VCC VCC _2039_
+ sky130_fd_sc_hs__and2b_1
X_5596_ clknet_leaf_36_i_clk _0243_ VSS VSS VCC VCC u_muldiv.mul\[13\] sky130_fd_sc_hs__dfxtp_1
X_4547_ _1214_ VSS VSS VCC VCC _2006_ sky130_fd_sc_hs__buf_2
X_4478_ u_muldiv.divisor\[62\] _1210_ _1970_ u_bits.i_op2\[31\] VSS VSS VCC
+ VCC _0228_ sky130_fd_sc_hs__a22o_1
X_3429_ op_cnt\[1\] _1197_ _1198_ VSS VSS VCC VCC _1199_ sky130_fd_sc_hs__or3b_1
Xclkbuf_leaf_20_i_clk clknet_2_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_20_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_2800_ _0496_ _0614_ VSS VSS VCC VCC _0615_ sky130_fd_sc_hs__nand2_2
X_3780_ _1110_ _1085_ _1500_ _1248_ _1502_ VSS VSS VCC VCC _1503_ sky130_fd_sc_hs__a221o_1
X_2731_ _0530_ _0531_ VSS VSS VCC VCC _0546_ sky130_fd_sc_hs__nand2_1
Xclkbuf_leaf_35_i_clk clknet_2_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_35_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5450_ clknet_leaf_9_i_clk _0098_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[10\]
+ sky130_fd_sc_hs__dfxtp_1
X_2662_ u_bits.i_op1\[18\] u_muldiv.add_prev\[18\] _0451_ VSS VSS VCC VCC
+ _0477_ sky130_fd_sc_hs__mux2_1
X_4401_ u_muldiv.divisor\[46\] _1867_ _1887_ u_muldiv.divisor\[47\] _1909_ VSS VSS
+ VCC VCC _0212_ sky130_fd_sc_hs__a221o_1
X_5381_ clknet_leaf_48_i_clk _0029_ VSS VSS VCC VCC u_bits.i_op1\[13\] sky130_fd_sc_hs__dfxtp_2
X_4332_ _1851_ _1853_ VSS VSS VCC VCC _1854_ sky130_fd_sc_hs__nor2_1
X_4263_ csr_data\[14\] i_csr_data[14] _1800_ VSS VSS VCC VCC _1806_ sky130_fd_sc_hs__mux2_1
X_3214_ _0987_ _0988_ VSS VSS VCC VCC _1014_ sky130_fd_sc_hs__nand2_1
X_4194_ _1770_ VSS VSS VCC VCC _0144_ sky130_fd_sc_hs__clkbuf_1
X_3145_ _0943_ u_bits.i_op2\[25\] VSS VSS VCC VCC _0950_ sky130_fd_sc_hs__nand2_1
X_3076_ _0858_ _0865_ _0869_ _0884_ VSS VSS VCC VCC _0885_ sky130_fd_sc_hs__or4_1
X_3978_ _1635_ VSS VSS VCC VCC _1641_ sky130_fd_sc_hs__buf_2
X_2929_ _0633_ VSS VSS VCC VCC _0742_ sky130_fd_sc_hs__buf_2
X_5717_ clknet_leaf_24_i_clk _0360_ VSS VSS VCC VCC u_muldiv.dividend\[1\]
+ sky130_fd_sc_hs__dfxtp_2
X_5648_ clknet_leaf_10_i_clk _0292_ VSS VSS VCC VCC op_cnt\[0\] sky130_fd_sc_hs__dfxtp_1
X_5579_ clknet_leaf_9_i_clk _0226_ VSS VSS VCC VCC u_muldiv.divisor\[60\]
+ sky130_fd_sc_hs__dfxtp_1
X_4950_ _2295_ _2308_ _1255_ VSS VSS VCC VCC _2310_ sky130_fd_sc_hs__a21oi_1
X_4881_ u_muldiv.o_div\[30\] _2274_ _2244_ VSS VSS VCC VCC _2275_ sky130_fd_sc_hs__mux2_1
X_3901_ _1310_ i_op1[4] _1599_ VSS VSS VCC VCC _1602_ sky130_fd_sc_hs__mux2_1
X_3832_ _1541_ _1551_ _0446_ VSS VSS VCC VCC _1552_ sky130_fd_sc_hs__a21o_1
X_5502_ clknet_leaf_43_i_clk _0150_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[20\]
+ sky130_fd_sc_hs__dfxtp_1
X_3763_ u_bits.i_op2\[13\] VSS VSS VCC VCC _1487_ sky130_fd_sc_hs__clkbuf_4
X_2714_ _0459_ u_bits.i_op2\[2\] u_bits.i_op1\[2\] _0463_ VSS VSS VCC VCC
+ _0529_ sky130_fd_sc_hs__a22o_1
X_3694_ u_bits.i_op2\[8\] _0785_ _1272_ VSS VSS VCC VCC _1423_ sky130_fd_sc_hs__a21oi_1
X_2645_ _0459_ VSS VSS VCC VCC _0460_ sky130_fd_sc_hs__buf_2
X_5433_ clknet_leaf_0_i_clk _0081_ VSS VSS VCC VCC u_bits.i_op2\[24\] sky130_fd_sc_hs__dfxtp_2
X_5364_ clknet_leaf_34_i_clk _0012_ VSS VSS VCC VCC u_muldiv.mul\[60\] sky130_fd_sc_hs__dfxtp_1
X_4315_ _1835_ VSS VSS VCC VCC _1838_ sky130_fd_sc_hs__buf_2
X_5295_ u_muldiv.divisor\[9\] _2614_ _2615_ u_muldiv.divisor\[10\] VSS VSS VCC
+ VCC _0400_ sky130_fd_sc_hs__a22o_1
X_4246_ csr_data\[6\] i_csr_data[6] _1789_ VSS VSS VCC VCC _1797_ sky130_fd_sc_hs__mux2_1
X_4177_ _1761_ VSS VSS VCC VCC _0136_ sky130_fd_sc_hs__clkbuf_1
X_3128_ _0458_ _0933_ VSS VSS VCC VCC _0934_ sky130_fd_sc_hs__xnor2_4
X_3059_ _0692_ u_bits.i_op2\[23\] _0867_ VSS VSS VCC VCC _0868_ sky130_fd_sc_hs__a21oi_1
X_5080_ _0776_ _2293_ _2428_ VSS VSS VCC VCC _2429_ sky130_fd_sc_hs__nand3_1
X_4100_ _1722_ VSS VSS VCC VCC _0098_ sky130_fd_sc_hs__clkbuf_1
X_4031_ _1665_ _1677_ _1678_ VSS VSS VCC VCC _0073_ sky130_fd_sc_hs__a21o_1
X_4933_ _0917_ _0791_ _2293_ u_muldiv.on_wait VSS VSS VCC VCC _2294_ sky130_fd_sc_hs__a31o_1
X_4864_ u_muldiv.quotient_msk\[27\] _2258_ _2229_ VSS VSS VCC VCC _2261_ sky130_fd_sc_hs__mux2_1
X_4795_ u_muldiv.quotient_msk\[13\] _2201_ _2156_ VSS VSS VCC VCC _2206_ sky130_fd_sc_hs__mux2_1
X_3815_ _0628_ _1529_ _1532_ _1535_ VSS VSS VCC VCC _1536_ sky130_fd_sc_hs__or4_1
X_3746_ _0788_ _1470_ VSS VSS VCC VCC _1471_ sky130_fd_sc_hs__or2_1
X_5416_ clknet_leaf_46_i_clk _0064_ VSS VSS VCC VCC u_bits.i_op2\[7\] sky130_fd_sc_hs__dfxtp_1
X_3677_ _1406_ _1258_ _0867_ VSS VSS VCC VCC _1407_ sky130_fd_sc_hs__a21oi_1
X_5347_ _1163_ _2628_ VSS VSS VCC VCC _0439_ sky130_fd_sc_hs__nor2_1
X_5278_ _2607_ _2608_ VSS VSS VCC VCC _2609_ sky130_fd_sc_hs__xnor2_1
X_4229_ _1788_ VSS VSS VCC VCC _0161_ sky130_fd_sc_hs__clkbuf_1
X_3600_ _1106_ csr_data\[2\] _1124_ VSS VSS VCC VCC _1335_ sky130_fd_sc_hs__o21ai_1
X_4580_ _2014_ VSS VSS VCC VCC _0286_ sky130_fd_sc_hs__clkbuf_1
X_3531_ _0831_ _0917_ _1267_ VSS VSS VCC VCC _1268_ sky130_fd_sc_hs__a21oi_1
X_3462_ _1221_ VSS VSS VCC VCC o_wdata[13] sky130_fd_sc_hs__buf_2
X_5201_ _0904_ _2293_ _2537_ VSS VSS VCC VCC _2539_ sky130_fd_sc_hs__and3_1
X_3393_ _1095_ _1099_ VSS VSS VCC VCC _1168_ sky130_fd_sc_hs__nand2_1
X_5132_ u_muldiv.dividend\[18\] _2468_ VSS VSS VCC VCC _2476_ sky130_fd_sc_hs__xor2_1
X_5063_ _2413_ VSS VSS VCC VCC _0370_ sky130_fd_sc_hs__clkbuf_1
X_4014_ u_bits.i_op2\[11\] _1663_ _1651_ i_op2[11] VSS VSS VCC VCC _1667_
+ sky130_fd_sc_hs__a22o_1
X_4916_ u_muldiv.quotient_msk\[24\] _2282_ _2283_ u_muldiv.quotient_msk\[25\] VSS
+ VSS VCC VCC _0353_ sky130_fd_sc_hs__a22o_1
X_4847_ _2161_ _2247_ u_muldiv.o_div\[23\] VSS VSS VCC VCC _2248_ sky130_fd_sc_hs__a21oi_1
X_4778_ _2181_ _2190_ _2192_ VSS VSS VCC VCC _0306_ sky130_fd_sc_hs__a21oi_1
X_3729_ _1333_ csr_data\[10\] _1388_ VSS VSS VCC VCC _1456_ sky130_fd_sc_hs__o21ai_1
X_5750_ clknet_leaf_24_i_clk _0393_ VSS VSS VCC VCC u_muldiv.divisor\[2\]
+ sky130_fd_sc_hs__dfxtp_1
X_2962_ _0772_ _0773_ _0774_ VSS VSS VCC VCC _0775_ sky130_fd_sc_hs__mux2_2
X_5681_ clknet_leaf_31_i_clk _0324_ VSS VSS VCC VCC u_muldiv.o_div\[27\] sky130_fd_sc_hs__dfxtp_1
X_4701_ _2123_ u_muldiv.dividend\[27\] u_muldiv.dividend\[26\] VSS VSS VCC VCC
+ _2124_ sky130_fd_sc_hs__o21ai_1
X_4632_ u_muldiv.dividend\[7\] u_muldiv.divisor\[7\] VSS VSS VCC VCC _2055_
+ sky130_fd_sc_hs__and2b_1
X_2893_ _0695_ _0706_ _0707_ VSS VSS VCC VCC _0708_ sky130_fd_sc_hs__mux2_1
X_4563_ o_add[16] _2004_ VSS VSS VCC VCC _2008_ sky130_fd_sc_hs__and2_1
X_4494_ _1583_ VSS VSS VCC VCC _1978_ sky130_fd_sc_hs__clkbuf_4
X_3514_ u_bits.i_op1\[11\] VSS VSS VCC VCC _1251_ sky130_fd_sc_hs__buf_4
X_3445_ _1204_ i_alu_ctrl[1] _1202_ _1211_ VSS VSS VCC VCC _1212_ sky130_fd_sc_hs__o2bb2a_1
X_3376_ _1153_ _1156_ VSS VSS VCC VCC _1157_ sky130_fd_sc_hs__nand2_4
X_5115_ _0653_ _2460_ VSS VSS VCC VCC _2461_ sky130_fd_sc_hs__xnor2_1
X_5046_ _2051_ _2077_ _2050_ VSS VSS VCC VCC _2398_ sky130_fd_sc_hs__o21ai_1
X_3230_ u_bits.i_op1\[28\] VSS VSS VCC VCC _1029_ sky130_fd_sc_hs__clkbuf_4
X_3161_ _0898_ _0899_ _0934_ _0935_ VSS VSS VCC VCC _0965_ sky130_fd_sc_hs__a22o_1
X_3092_ _0898_ _0899_ VSS VSS VCC VCC _0900_ sky130_fd_sc_hs__xnor2_1
X_5802_ clknet_leaf_39_i_clk _0444_ VSS VSS VCC VCC u_muldiv.mul\[50\] sky130_fd_sc_hs__dfxtp_1
X_3994_ _1641_ _1650_ _1652_ VSS VSS VCC VCC _0062_ sky130_fd_sc_hs__a21o_1
X_5733_ clknet_leaf_18_i_clk _0376_ VSS VSS VCC VCC u_muldiv.dividend\[17\]
+ sky130_fd_sc_hs__dfxtp_2
X_2945_ u_bits.i_op2\[2\] VSS VSS VCC VCC _0758_ sky130_fd_sc_hs__clkbuf_4
X_5664_ clknet_leaf_28_i_clk _0307_ VSS VSS VCC VCC u_muldiv.o_div\[10\] sky130_fd_sc_hs__dfxtp_1
X_2876_ u_bits.i_op1\[22\] VSS VSS VCC VCC _0691_ sky130_fd_sc_hs__buf_4
X_4615_ u_muldiv.divisor\[18\] _2037_ u_muldiv.dividend\[18\] VSS VSS VCC VCC
+ _2038_ sky130_fd_sc_hs__or3b_1
X_5595_ clknet_leaf_36_i_clk _0242_ VSS VSS VCC VCC u_muldiv.mul\[12\] sky130_fd_sc_hs__dfxtp_1
X_4546_ _2005_ VSS VSS VCC VCC _0261_ sky130_fd_sc_hs__clkbuf_1
X_4477_ _1868_ _1969_ _1833_ VSS VSS VCC VCC _1970_ sky130_fd_sc_hs__a21oi_1
X_3428_ u_muldiv.i_is_div VSS VSS VCC VCC _1198_ sky130_fd_sc_hs__buf_4
X_3359_ _0594_ _1144_ VSS VSS VCC VCC _1145_ sky130_fd_sc_hs__xor2_4
X_5029_ _2052_ _2371_ VSS VSS VCC VCC _2382_ sky130_fd_sc_hs__nand2_1
Xclkbuf_2_1__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_1__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
Xclkbuf_leaf_1_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_1_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_2730_ _0526_ _0527_ VSS VSS VCC VCC _0545_ sky130_fd_sc_hs__nand2_1
X_2661_ _0457_ _0475_ VSS VSS VCC VCC _0476_ sky130_fd_sc_hs__xnor2_1
X_4400_ _1907_ _1908_ VSS VSS VCC VCC _1909_ sky130_fd_sc_hs__nor2_1
X_5380_ clknet_leaf_48_i_clk _0028_ VSS VSS VCC VCC u_bits.i_op1\[12\] sky130_fd_sc_hs__dfxtp_2
X_4331_ _0923_ _0915_ _1852_ _1832_ VSS VSS VCC VCC _1853_ sky130_fd_sc_hs__a31o_1
X_4262_ _1805_ VSS VSS VCC VCC _0177_ sky130_fd_sc_hs__clkbuf_1
X_3213_ _0964_ _0991_ VSS VSS VCC VCC _1013_ sky130_fd_sc_hs__nand2_1
X_4193_ u_wr_mux.i_reg_data2\[14\] i_reg_data2[14] _1767_ VSS VSS VCC VCC
+ _1770_ sky130_fd_sc_hs__mux2_1
X_3144_ _0947_ _0948_ _0707_ VSS VSS VCC VCC _0949_ sky130_fd_sc_hs__mux2_1
X_3075_ _0643_ _0878_ _0883_ _0800_ VSS VSS VCC VCC _0884_ sky130_fd_sc_hs__o211a_1
X_3977_ _0831_ _1637_ _1638_ i_op2[0] _1640_ VSS VSS VCC VCC _0057_ sky130_fd_sc_hs__a221o_1
X_5716_ clknet_leaf_36_i_clk _0359_ VSS VSS VCC VCC u_muldiv.quotient_msk\[30\]
+ sky130_fd_sc_hs__dfxtp_1
X_2928_ _0719_ VSS VSS VCC VCC _0741_ sky130_fd_sc_hs__buf_2
X_5647_ clknet_leaf_8_i_clk _0000_ VSS VSS VCC VCC u_muldiv.i_on_end sky130_fd_sc_hs__dfxtp_2
X_2859_ _0673_ VSS VSS VCC VCC _0674_ sky130_fd_sc_hs__clkbuf_4
X_5578_ clknet_leaf_9_i_clk _0225_ VSS VSS VCC VCC u_muldiv.divisor\[59\]
+ sky130_fd_sc_hs__dfxtp_1
X_4529_ _1996_ VSS VSS VCC VCC _0253_ sky130_fd_sc_hs__clkbuf_1
X_4880_ _2271_ _2272_ _2273_ _1841_ VSS VSS VCC VCC _2274_ sky130_fd_sc_hs__a22o_1
X_3900_ _1601_ VSS VSS VCC VCC _0019_ sky130_fd_sc_hs__clkbuf_1
X_3831_ _0749_ o_add[17] _1549_ _1550_ _0453_ VSS VSS VCC VCC _1551_ sky130_fd_sc_hs__a221o_1
X_3762_ _0759_ _1485_ _0824_ _0765_ _0920_ _0643_ VSS VSS VCC VCC _1486_ sky130_fd_sc_hs__mux4_1
X_5501_ clknet_leaf_43_i_clk _0149_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[19\]
+ sky130_fd_sc_hs__dfxtp_1
X_2713_ _0526_ _0527_ VSS VSS VCC VCC _0528_ sky130_fd_sc_hs__nor2_1
X_3693_ _0908_ _1421_ VSS VSS VCC VCC _1422_ sky130_fd_sc_hs__nor2_1
X_2644_ u_mux.i_group_mux VSS VSS VCC VCC _0459_ sky130_fd_sc_hs__inv_2
X_5432_ clknet_leaf_0_i_clk _0080_ VSS VSS VCC VCC u_bits.i_op2\[23\] sky130_fd_sc_hs__dfxtp_4
X_5363_ clknet_leaf_39_i_clk _0011_ VSS VSS VCC VCC u_muldiv.mul\[59\] sky130_fd_sc_hs__dfxtp_1
X_4314_ u_muldiv.divisor\[32\] _1829_ _1833_ _0831_ _1837_ VSS VSS VCC VCC
+ _0197_ sky130_fd_sc_hs__o221a_1
X_5294_ _1842_ VSS VSS VCC VCC _2615_ sky130_fd_sc_hs__buf_2
X_4245_ _1796_ VSS VSS VCC VCC _0169_ sky130_fd_sc_hs__clkbuf_1
X_4176_ o_wdata[6] i_reg_data2[6] _1756_ VSS VSS VCC VCC _1761_ sky130_fd_sc_hs__mux2_1
X_3127_ _0461_ u_bits.i_op2\[25\] _0465_ u_bits.i_op1\[25\] VSS VSS VCC VCC
+ _0933_ sky130_fd_sc_hs__a22o_1
X_3058_ _0866_ VSS VSS VCC VCC _0867_ sky130_fd_sc_hs__buf_2
Xclkbuf_leaf_34_i_clk clknet_2_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_34_i_clk
+ sky130_fd_sc_hs__clkbuf_16
Xclkbuf_leaf_49_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_49_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4030_ u_bits.i_op2\[16\] _1663_ _1675_ i_op2[16] VSS VSS VCC VCC _1678_
+ sky130_fd_sc_hs__a22o_1
X_4932_ _2292_ VSS VSS VCC VCC _2293_ sky130_fd_sc_hs__buf_2
X_4863_ u_muldiv.o_div\[27\] _2170_ _2258_ _2196_ VSS VSS VCC VCC _2260_ sky130_fd_sc_hs__a31o_1
X_4794_ _2170_ u_muldiv.o_div\[13\] _2201_ _2196_ VSS VSS VCC VCC _2205_ sky130_fd_sc_hs__a31o_1
X_3814_ _0672_ _1533_ _1534_ _0800_ VSS VSS VCC VCC _1535_ sky130_fd_sc_hs__o211a_1
X_3745_ _1253_ _1261_ _0668_ VSS VSS VCC VCC _1470_ sky130_fd_sc_hs__mux2_1
X_3676_ u_bits.i_op2\[7\] VSS VSS VCC VCC _1406_ sky130_fd_sc_hs__buf_4
X_5415_ clknet_leaf_49_i_clk _0063_ VSS VSS VCC VCC u_bits.i_op2\[6\] sky130_fd_sc_hs__dfxtp_4
X_5346_ _1155_ _2628_ VSS VSS VCC VCC _0438_ sky130_fd_sc_hs__nor2_1
X_5277_ _2137_ _2144_ VSS VSS VCC VCC _2608_ sky130_fd_sc_hs__nor2_1
X_4228_ u_wr_mux.i_reg_data2\[31\] i_reg_data2[31] _1778_ VSS VSS VCC VCC
+ _1788_ sky130_fd_sc_hs__mux2_1
X_4159_ u_bits.i_sra i_alu_ctrl[3] _1745_ VSS VSS VCC VCC _1752_ sky130_fd_sc_hs__mux2_1
X_3530_ _0867_ VSS VSS VCC VCC _1267_ sky130_fd_sc_hs__clkbuf_4
X_3461_ u_wr_mux.i_reg_data2\[13\] o_wdata[5] _0718_ VSS VSS VCC VCC _1221_
+ sky130_fd_sc_hs__mux2_1
X_5200_ _2295_ _2537_ _0904_ VSS VSS VCC VCC _2538_ sky130_fd_sc_hs__a21oi_1
X_3392_ _1095_ _1099_ VSS VSS VCC VCC _1167_ sky130_fd_sc_hs__nor2_1
X_5131_ _2475_ VSS VSS VCC VCC _0376_ sky130_fd_sc_hs__clkbuf_1
X_5062_ u_muldiv.dividend\[11\] _2412_ _2378_ VSS VSS VCC VCC _2413_ sky130_fd_sc_hs__mux2_1
X_4013_ u_bits.i_op2\[12\] _1445_ _1657_ VSS VSS VCC VCC _1666_ sky130_fd_sc_hs__mux2_1
X_4915_ u_muldiv.quotient_msk\[23\] _2282_ _2283_ u_muldiv.quotient_msk\[24\] VSS
+ VSS VCC VCC _0352_ sky130_fd_sc_hs__a22o_1
X_4846_ u_muldiv.quotient_msk\[23\] _2241_ _2229_ VSS VSS VCC VCC _2247_ sky130_fd_sc_hs__mux2_1
X_4777_ _2167_ _2191_ u_muldiv.o_div\[9\] VSS VSS VCC VCC _2192_ sky130_fd_sc_hs__a21oi_1
X_3728_ _1331_ _1451_ _1453_ _1454_ _1357_ VSS VSS VCC VCC _1455_ sky130_fd_sc_hs__o221a_1
X_3659_ _1309_ _1314_ _1312_ _1306_ _0669_ _0920_ VSS VSS VCC VCC _1390_ sky130_fd_sc_hs__mux4_1
X_5329_ _2625_ VSS VSS VCC VCC _0424_ sky130_fd_sc_hs__clkbuf_1
X_2961_ _0659_ VSS VSS VCC VCC _0774_ sky130_fd_sc_hs__clkbuf_4
X_5680_ clknet_leaf_31_i_clk _0323_ VSS VSS VCC VCC u_muldiv.o_div\[26\] sky130_fd_sc_hs__dfxtp_1
X_4700_ u_muldiv.divisor\[27\] VSS VSS VCC VCC _2123_ sky130_fd_sc_hs__inv_2
X_4631_ _2052_ _2053_ VSS VSS VCC VCC _2054_ sky130_fd_sc_hs__nand2_1
X_2892_ _0524_ VSS VSS VCC VCC _0707_ sky130_fd_sc_hs__clkbuf_4
X_4562_ _1162_ _2007_ VSS VSS VCC VCC _0275_ sky130_fd_sc_hs__nor2_1
X_4493_ _1977_ VSS VSS VCC VCC _0236_ sky130_fd_sc_hs__clkbuf_1
X_3513_ u_bits.i_op1\[9\] VSS VSS VCC VCC _1250_ sky130_fd_sc_hs__buf_4
X_3444_ u_muldiv.i_on_wait VSS VSS VCC VCC _1211_ sky130_fd_sc_hs__clkinv_2
X_3375_ _0578_ _1152_ _0607_ VSS VSS VCC VCC _1156_ sky130_fd_sc_hs__nand3_1
X_5114_ _0654_ _2450_ _2385_ VSS VSS VCC VCC _2460_ sky130_fd_sc_hs__o21ai_1
X_5045_ _2050_ _2051_ _2077_ VSS VSS VCC VCC _2397_ sky130_fd_sc_hs__or3_1
X_4829_ u_muldiv.o_div\[20\] u_muldiv.o_div\[19\] _2226_ VSS VSS VCC VCC _2233_
+ sky130_fd_sc_hs__or3_2
X_3160_ _0962_ _0963_ VSS VSS VCC VCC _0964_ sky130_fd_sc_hs__and2_2
X_3091_ u_bits.i_op1\[24\] u_muldiv.add_prev\[24\] _0452_ VSS VSS VCC VCC
+ _0899_ sky130_fd_sc_hs__mux2_1
X_5801_ clknet_leaf_35_i_clk _0443_ VSS VSS VCC VCC u_muldiv.mul\[49\] sky130_fd_sc_hs__dfxtp_1
X_5732_ clknet_leaf_18_i_clk _0375_ VSS VSS VCC VCC u_muldiv.dividend\[16\]
+ sky130_fd_sc_hs__dfxtp_2
X_3993_ _1376_ _1637_ _1651_ i_op2[5] VSS VSS VCC VCC _1652_ sky130_fd_sc_hs__a22o_1
X_2944_ _0755_ _0756_ _0648_ VSS VSS VCC VCC _0757_ sky130_fd_sc_hs__mux2_1
X_5663_ clknet_leaf_27_i_clk _0306_ VSS VSS VCC VCC u_muldiv.o_div\[9\] sky130_fd_sc_hs__dfxtp_1
X_2875_ u_bits.i_op1\[24\] u_bits.i_op1\[25\] _0689_ u_bits.i_op1\[27\] _0650_ _0659_
+ VSS VSS VCC VCC _0690_ sky130_fd_sc_hs__mux4_1
X_4614_ u_muldiv.dividend\[19\] u_muldiv.divisor\[19\] VSS VSS VCC VCC _2037_
+ sky130_fd_sc_hs__and2b_1
X_5594_ clknet_leaf_36_i_clk _0241_ VSS VSS VCC VCC u_muldiv.mul\[11\] sky130_fd_sc_hs__dfxtp_1
X_4545_ o_add[1] _2004_ VSS VSS VCC VCC _2005_ sky130_fd_sc_hs__and2_1
X_4476_ u_bits.i_op2\[29\] u_bits.i_op2\[30\] _1962_ VSS VSS VCC VCC _1969_
+ sky130_fd_sc_hs__or3_1
X_3427_ op_cnt\[2\] op_cnt\[3\] op_cnt\[4\] op_cnt\[5\] VSS VSS VCC VCC _1197_
+ sky130_fd_sc_hs__or4b_1
X_3358_ _0596_ _0597_ _1143_ VSS VSS VCC VCC _1144_ sky130_fd_sc_hs__a21bo_1
X_3289_ _0832_ _0833_ _1083_ _0976_ _0825_ _0920_ VSS VSS VCC VCC _1084_ sky130_fd_sc_hs__mux4_1
X_5028_ u_muldiv.dividend\[8\] _2361_ u_muldiv.dividend\[9\] VSS VSS VCC VCC
+ _2381_ sky130_fd_sc_hs__o21ai_1
X_2660_ _0460_ u_bits.i_op2\[18\] u_bits.i_op1\[18\] _0464_ VSS VSS VCC VCC
+ _0475_ sky130_fd_sc_hs__a22o_1
X_4330_ _1845_ VSS VSS VCC VCC _1852_ sky130_fd_sc_hs__buf_2
X_4261_ csr_data\[13\] i_csr_data[13] _1800_ VSS VSS VCC VCC _1805_ sky130_fd_sc_hs__mux2_1
X_3212_ _0739_ csr_data\[27\] _1012_ _0732_ VSS VSS VCC VCC o_result[27] sky130_fd_sc_hs__o211a_2
X_4192_ _1769_ VSS VSS VCC VCC _0143_ sky130_fd_sc_hs__clkbuf_1
X_3143_ _0669_ _0793_ VSS VSS VCC VCC _0948_ sky130_fd_sc_hs__nor2_1
X_3074_ _0879_ _0882_ _0642_ VSS VSS VCC VCC _0883_ sky130_fd_sc_hs__a21bo_1
X_3976_ _1639_ _1635_ _1112_ VSS VSS VCC VCC _1640_ sky130_fd_sc_hs__and3b_1
X_5715_ clknet_leaf_32_i_clk _0358_ VSS VSS VCC VCC u_muldiv.quotient_msk\[29\]
+ sky130_fd_sc_hs__dfxtp_1
X_2927_ _0622_ VSS VSS VCC VCC _0740_ sky130_fd_sc_hs__buf_2
X_5646_ clknet_leaf_11_i_clk _0002_ VSS VSS VCC VCC u_muldiv.i_on_wait sky130_fd_sc_hs__dfxtp_2
X_2858_ _0524_ VSS VSS VCC VCC _0673_ sky130_fd_sc_hs__inv_2
X_5577_ clknet_leaf_9_i_clk _0224_ VSS VSS VCC VCC u_muldiv.divisor\[58\]
+ sky130_fd_sc_hs__dfxtp_1
X_2789_ _0592_ _0593_ _0596_ _0597_ VSS VSS VCC VCC _0604_ sky130_fd_sc_hs__a22o_1
X_4528_ u_muldiv.mul\[23\] u_muldiv.mul\[24\] _1989_ VSS VSS VCC VCC _1996_
+ sky130_fd_sc_hs__mux2_1
X_4459_ u_bits.i_op2\[27\] _1955_ _1832_ VSS VSS VCC VCC _1956_ sky130_fd_sc_hs__a21oi_1
X_3830_ _0629_ _1543_ _0955_ VSS VSS VCC VCC _1550_ sky130_fd_sc_hs__a21oi_1
X_3761_ _1282_ _1288_ _0758_ VSS VSS VCC VCC _1485_ sky130_fd_sc_hs__mux2_1
X_2712_ u_bits.i_op1\[3\] u_muldiv.add_prev\[3\] _0450_ VSS VSS VCC VCC _0527_
+ sky130_fd_sc_hs__mux2_1
X_5500_ clknet_leaf_43_i_clk _0148_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[18\]
+ sky130_fd_sc_hs__dfxtp_1
X_3692_ _1110_ _0921_ _1418_ _1249_ _1420_ VSS VSS VCC VCC _1421_ sky130_fd_sc_hs__a221o_1
X_2643_ _0457_ VSS VSS VCC VCC _0458_ sky130_fd_sc_hs__buf_4
X_5431_ clknet_leaf_0_i_clk _0079_ VSS VSS VCC VCC u_bits.i_op2\[22\] sky130_fd_sc_hs__dfxtp_4
X_5362_ clknet_leaf_40_i_clk _0010_ VSS VSS VCC VCC u_muldiv.mul\[58\] sky130_fd_sc_hs__dfxtp_1
X_4313_ _1834_ _1836_ VSS VSS VCC VCC _1837_ sky130_fd_sc_hs__nand2_1
X_5293_ u_muldiv.divisor\[8\] _2614_ _2285_ u_muldiv.divisor\[9\] VSS VSS VCC
+ VCC _0399_ sky130_fd_sc_hs__a22o_1
Xclkbuf_leaf_0_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_0_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4244_ csr_data\[5\] i_csr_data[5] _1789_ VSS VSS VCC VCC _1796_ sky130_fd_sc_hs__mux2_1
X_4175_ _1760_ VSS VSS VCC VCC _0135_ sky130_fd_sc_hs__clkbuf_1
X_3126_ _0739_ csr_data\[24\] _0932_ _0732_ VSS VSS VCC VCC o_result[24] sky130_fd_sc_hs__o211a_2
X_3057_ o_funct3[2] _0638_ VSS VSS VCC VCC _0866_ sky130_fd_sc_hs__nand2_1
X_3959_ _1596_ VSS VSS VCC VCC _1632_ sky130_fd_sc_hs__clkbuf_4
X_5629_ clknet_leaf_44_i_clk _0276_ VSS VSS VCC VCC u_muldiv.add_prev\[15\]
+ sky130_fd_sc_hs__dfxtp_1
X_4931_ _2291_ VSS VSS VCC VCC _2292_ sky130_fd_sc_hs__buf_2
X_4862_ u_muldiv.o_div\[26\] _2171_ _2259_ _2164_ VSS VSS VCC VCC _0323_ sky130_fd_sc_hs__a22o_1
X_3813_ _0672_ _1266_ VSS VSS VCC VCC _1534_ sky130_fd_sc_hs__nand2_1
X_4793_ _2204_ VSS VSS VCC VCC _0309_ sky130_fd_sc_hs__clkbuf_1
X_3744_ _1468_ _1469_ _1336_ u_pc_sel.i_pc_next\[11\] VSS VSS VCC VCC o_result[11]
+ sky130_fd_sc_hs__a2bb2o_2
X_3675_ _1404_ _0864_ _0751_ VSS VSS VCC VCC _1405_ sky130_fd_sc_hs__mux2_1
X_5414_ clknet_leaf_49_i_clk _0062_ VSS VSS VCC VCC u_bits.i_op2\[5\] sky130_fd_sc_hs__dfxtp_1
X_5345_ _1157_ _2628_ VSS VSS VCC VCC _0437_ sky130_fd_sc_hs__nor2_1
X_5276_ _2136_ u_muldiv.dividend\[30\] _2135_ VSS VSS VCC VCC _2607_ sky130_fd_sc_hs__a21oi_1
X_4227_ _1787_ VSS VSS VCC VCC _0160_ sky130_fd_sc_hs__clkbuf_1
X_4158_ _1751_ VSS VSS VCC VCC _0127_ sky130_fd_sc_hs__clkbuf_1
X_3109_ u_bits.i_op2\[2\] _0915_ VSS VSS VCC VCC _0916_ sky130_fd_sc_hs__or2_2
X_4089_ u_pc_sel.i_pc_next\[5\] i_pc_next[5] _1712_ VSS VSS VCC VCC _1717_
+ sky130_fd_sc_hs__mux2_1
X_3460_ _1220_ VSS VSS VCC VCC o_wdata[12] sky130_fd_sc_hs__buf_2
X_3391_ _0616_ VSS VSS VCC VCC o_add[20] sky130_fd_sc_hs__inv_2
X_5130_ u_muldiv.dividend\[17\] _2474_ _2378_ VSS VSS VCC VCC _2475_ sky130_fd_sc_hs__mux2_1
X_5061_ _1208_ _2403_ _2404_ _2408_ _2411_ VSS VSS VCC VCC _2412_ sky130_fd_sc_hs__a32o_1
X_4012_ _1635_ VSS VSS VCC VCC _1665_ sky130_fd_sc_hs__buf_2
X_4914_ u_muldiv.quotient_msk\[22\] _2282_ _2283_ u_muldiv.quotient_msk\[23\] VSS
+ VSS VCC VCC _0351_ sky130_fd_sc_hs__a22o_1
X_4845_ u_muldiv.o_div\[23\] _2170_ _2241_ _2196_ VSS VSS VCC VCC _2246_ sky130_fd_sc_hs__a31o_1
X_4776_ u_muldiv.quotient_msk\[9\] _2186_ _2156_ VSS VSS VCC VCC _2191_ sky130_fd_sc_hs__mux2_1
X_3727_ u_muldiv.mul\[10\] _1330_ _1400_ VSS VSS VCC VCC _1454_ sky130_fd_sc_hs__o21ai_1
Xclkbuf_leaf_33_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_33_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3658_ _1387_ _1389_ _1336_ u_pc_sel.i_pc_next\[5\] VSS VSS VCC VCC o_result[5]
+ sky130_fd_sc_hs__a2bb2o_2
X_3589_ _1274_ _1322_ _1323_ _0624_ _1130_ VSS VSS VCC VCC _1324_ sky130_fd_sc_hs__o32a_1
X_5328_ u_muldiv.dividend\[0\] _2624_ _2152_ VSS VSS VCC VCC _2625_ sky130_fd_sc_hs__mux2_1
Xclkbuf_leaf_48_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_48_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5259_ _1208_ _2583_ _2584_ _2591_ VSS VSS VCC VCC _2592_ sky130_fd_sc_hs__a31o_1
X_2960_ u_bits.i_op1\[19\] _0645_ _0656_ VSS VSS VCC VCC _0773_ sky130_fd_sc_hs__mux2_1
X_2891_ _0705_ VSS VSS VCC VCC _0706_ sky130_fd_sc_hs__clkinv_2
X_4630_ u_muldiv.dividend\[8\] u_muldiv.divisor\[8\] VSS VSS VCC VCC _2053_
+ sky130_fd_sc_hs__or2b_1
X_4561_ _1163_ _2007_ VSS VSS VCC VCC _0274_ sky130_fd_sc_hs__nor2_1
X_4492_ u_muldiv.mul\[6\] u_muldiv.mul\[7\] _1584_ VSS VSS VCC VCC _1977_
+ sky130_fd_sc_hs__mux2_1
X_3512_ _1248_ VSS VSS VCC VCC _1249_ sky130_fd_sc_hs__clkbuf_4
X_3443_ _1204_ _1205_ _1210_ i_flush VSS VSS VCC VCC _0001_ sky130_fd_sc_hs__a211o_1
X_5113_ _2458_ _2089_ VSS VSS VCC VCC _2459_ sky130_fd_sc_hs__xor2_1
X_3374_ _1155_ VSS VSS VCC VCC o_add[13] sky130_fd_sc_hs__inv_2
X_5044_ _2295_ _2394_ _1305_ VSS VSS VCC VCC _2396_ sky130_fd_sc_hs__a21o_1
X_4828_ u_muldiv.o_div\[19\] _2226_ u_muldiv.o_div\[20\] VSS VSS VCC VCC _2232_
+ sky130_fd_sc_hs__o21ai_1
X_4759_ _2164_ _2175_ _2177_ VSS VSS VCC VCC _0302_ sky130_fd_sc_hs__a21oi_1
X_3090_ _0458_ _0897_ VSS VSS VCC VCC _0898_ sky130_fd_sc_hs__xnor2_2
X_3992_ _1595_ VSS VSS VCC VCC _1651_ sky130_fd_sc_hs__buf_2
X_5800_ clknet_leaf_39_i_clk _0442_ VSS VSS VCC VCC u_muldiv.mul\[48\] sky130_fd_sc_hs__dfxtp_1
X_5731_ clknet_leaf_21_i_clk _0374_ VSS VSS VCC VCC u_muldiv.dividend\[15\]
+ sky130_fd_sc_hs__dfxtp_2
X_2943_ u_bits.i_op1\[27\] u_bits.i_op1\[28\] _0649_ VSS VSS VCC VCC _0756_
+ sky130_fd_sc_hs__mux2_1
X_5662_ clknet_leaf_26_i_clk _0305_ VSS VSS VCC VCC u_muldiv.o_div\[8\] sky130_fd_sc_hs__dfxtp_1
X_2874_ u_bits.i_op1\[26\] VSS VSS VCC VCC _0689_ sky130_fd_sc_hs__buf_4
X_4613_ u_muldiv.divisor\[19\] u_muldiv.dividend\[19\] VSS VSS VCC VCC _2036_
+ sky130_fd_sc_hs__or2b_1
X_5593_ clknet_leaf_36_i_clk _0240_ VSS VSS VCC VCC u_muldiv.mul\[10\] sky130_fd_sc_hs__dfxtp_1
X_4544_ _1583_ VSS VSS VCC VCC _2004_ sky130_fd_sc_hs__clkbuf_4
X_4475_ u_muldiv.divisor\[61\] _1836_ _1946_ u_muldiv.divisor\[62\] _1968_ VSS VSS
+ VCC VCC _0227_ sky130_fd_sc_hs__a221o_1
X_3426_ u_pc_sel.i_inst_branch _1191_ _1196_ u_pc_sel.i_inst_jal_jalr VSS VSS
+ VCC VCC o_pc_select sky130_fd_sc_hs__a31o_2
X_3357_ _0568_ _0576_ _0598_ VSS VSS VCC VCC _1143_ sky130_fd_sc_hs__a21o_1
X_5027_ u_muldiv.dividend\[9\] u_muldiv.dividend\[8\] _2361_ VSS VSS VCC VCC
+ _2380_ sky130_fd_sc_hs__or3_1
X_3288_ _0699_ _0697_ _1029_ _0996_ _0651_ _0774_ VSS VSS VCC VCC _1083_ sky130_fd_sc_hs__mux4_1
X_4260_ _1804_ VSS VSS VCC VCC _0176_ sky130_fd_sc_hs__clkbuf_1
X_3211_ _0995_ _1011_ _0447_ VSS VSS VCC VCC _1012_ sky130_fd_sc_hs__a21o_1
X_4191_ u_wr_mux.i_reg_data2\[13\] i_reg_data2[13] _1767_ VSS VSS VCC VCC
+ _1769_ sky130_fd_sc_hs__mux2_1
X_3142_ _0787_ _0795_ _0758_ VSS VSS VCC VCC _0947_ sky130_fd_sc_hs__mux2_1
X_3073_ _0880_ _0881_ _0696_ VSS VSS VCC VCC _0882_ sky130_fd_sc_hs__mux2_1
X_3975_ _1198_ VSS VSS VCC VCC _1639_ sky130_fd_sc_hs__clkbuf_4
X_5714_ clknet_leaf_33_i_clk _0357_ VSS VSS VCC VCC u_muldiv.quotient_msk\[28\]
+ sky130_fd_sc_hs__dfxtp_1
X_2926_ _0728_ VSS VSS VCC VCC _0739_ sky130_fd_sc_hs__buf_2
X_5645_ clknet_leaf_9_i_clk _0001_ VSS VSS VCC VCC o_ready sky130_fd_sc_hs__dfxtp_2
X_2857_ _0642_ VSS VSS VCC VCC _0672_ sky130_fd_sc_hs__buf_2
X_5576_ clknet_leaf_9_i_clk _0223_ VSS VSS VCC VCC u_muldiv.divisor\[57\]
+ sky130_fd_sc_hs__dfxtp_1
X_2788_ _0587_ _0588_ VSS VSS VCC VCC _0603_ sky130_fd_sc_hs__nand2_1
X_4527_ _1995_ VSS VSS VCC VCC _0252_ sky130_fd_sc_hs__clkbuf_1
X_4458_ u_bits.i_op2\[26\] _1942_ _1951_ _1845_ VSS VSS VCC VCC _1955_ sky130_fd_sc_hs__o31a_1
X_3409_ _1135_ _1142_ _1147_ _1179_ VSS VSS VCC VCC _1180_ sky130_fd_sc_hs__and4_1
X_4389_ _1868_ _1899_ _1487_ VSS VSS VCC VCC _1900_ sky130_fd_sc_hs__a21oi_1
X_3760_ _1483_ _1484_ _0730_ u_pc_sel.i_pc_next\[12\] VSS VSS VCC VCC o_result[12]
+ sky130_fd_sc_hs__a2bb2o_2
X_2711_ _0457_ _0525_ VSS VSS VCC VCC _0526_ sky130_fd_sc_hs__xnor2_1
X_5430_ clknet_leaf_1_i_clk _0078_ VSS VSS VCC VCC u_bits.i_op2\[21\] sky130_fd_sc_hs__dfxtp_4
X_3691_ u_bits.i_op2\[8\] _0785_ _0637_ _1419_ VSS VSS VCC VCC _1420_ sky130_fd_sc_hs__o22a_1
X_2642_ _0456_ VSS VSS VCC VCC _0457_ sky130_fd_sc_hs__buf_4
X_5361_ clknet_leaf_39_i_clk _0009_ VSS VSS VCC VCC u_muldiv.mul\[57\] sky130_fd_sc_hs__dfxtp_1
X_5292_ u_muldiv.divisor\[7\] _2614_ _2285_ u_muldiv.divisor\[8\] VSS VSS VCC
+ VCC _0398_ sky130_fd_sc_hs__a22o_1
X_4312_ _1835_ VSS VSS VCC VCC _1836_ sky130_fd_sc_hs__buf_2
X_4243_ _1795_ VSS VSS VCC VCC _0168_ sky130_fd_sc_hs__clkbuf_1
X_4174_ o_wdata[5] i_reg_data2[5] _1756_ VSS VSS VCC VCC _1760_ sky130_fd_sc_hs__mux2_1
X_3125_ _0892_ _0931_ _0447_ VSS VSS VCC VCC _0932_ sky130_fd_sc_hs__a21o_1
X_3056_ _0643_ _0864_ _0711_ VSS VSS VCC VCC _0865_ sky130_fd_sc_hs__o21a_1
X_3958_ _1631_ VSS VSS VCC VCC _0047_ sky130_fd_sc_hs__clkbuf_1
X_3889_ i_flush i_reset_n o_ready VSS VSS VCC VCC _1594_ sky130_fd_sc_hs__and3b_1
X_2909_ _0461_ VSS VSS VCC VCC _0724_ sky130_fd_sc_hs__clkbuf_4
X_5628_ clknet_leaf_44_i_clk _0275_ VSS VSS VCC VCC u_muldiv.add_prev\[14\]
+ sky130_fd_sc_hs__dfxtp_1
X_5559_ clknet_leaf_7_i_clk _0206_ VSS VSS VCC VCC u_muldiv.divisor\[40\]
+ sky130_fd_sc_hs__dfxtp_1
X_4930_ _0620_ _0702_ VSS VSS VCC VCC _2291_ sky130_fd_sc_hs__and2b_1
X_4861_ _2165_ _2257_ _2258_ _1842_ u_muldiv.quotient_msk\[26\] VSS VSS VCC
+ VCC _2259_ sky130_fd_sc_hs__a32o_1
X_3812_ _0660_ _0664_ _0667_ _0678_ _0825_ _0707_ VSS VSS VCC VCC _1533_ sky130_fd_sc_hs__mux4_1
X_4792_ u_muldiv.o_div\[12\] _2203_ _2154_ VSS VSS VCC VCC _2204_ sky130_fd_sc_hs__mux2_1
X_3743_ _1333_ csr_data\[11\] _1388_ VSS VSS VCC VCC _1469_ sky130_fd_sc_hs__o21ai_1
X_3674_ _1339_ _1343_ _1341_ _1337_ _0669_ _0920_ VSS VSS VCC VCC _1404_ sky130_fd_sc_hs__mux4_1
X_5413_ clknet_leaf_49_i_clk _0061_ VSS VSS VCC VCC u_bits.i_op2\[4\] sky130_fd_sc_hs__dfxtp_2
X_5344_ _1150_ _2628_ VSS VSS VCC VCC _0436_ sky130_fd_sc_hs__nor2_1
X_5275_ u_muldiv.dividend\[31\] _2601_ _2605_ VSS VSS VCC VCC _2606_ sky130_fd_sc_hs__a21o_1
X_4226_ u_wr_mux.i_reg_data2\[30\] i_reg_data2[30] _1778_ VSS VSS VCC VCC
+ _1787_ sky130_fd_sc_hs__mux2_1
X_4157_ alu_ctrl\[2\] i_alu_ctrl[2] _1745_ VSS VSS VCC VCC _1751_ sky130_fd_sc_hs__mux2_1
X_3108_ u_bits.i_op2\[0\] u_bits.i_op2\[1\] VSS VSS VCC VCC _0915_ sky130_fd_sc_hs__or2_1
X_4088_ _1716_ VSS VSS VCC VCC _0092_ sky130_fd_sc_hs__clkbuf_1
X_3039_ _0458_ _0848_ VSS VSS VCC VCC _0849_ sky130_fd_sc_hs__xnor2_1
X_3390_ _0483_ _1165_ VSS VSS VCC VCC o_add[18] sky130_fd_sc_hs__xnor2_4
X_5060_ _2375_ _2410_ _1207_ VSS VSS VCC VCC _2411_ sky130_fd_sc_hs__a21oi_1
X_4011_ _1641_ _1662_ _1664_ VSS VSS VCC VCC _0067_ sky130_fd_sc_hs__a21o_1
X_4913_ u_muldiv.quotient_msk\[21\] _2282_ _2283_ u_muldiv.quotient_msk\[22\] VSS
+ VSS VCC VCC _0350_ sky130_fd_sc_hs__a22o_1
X_4844_ _2245_ VSS VSS VCC VCC _0319_ sky130_fd_sc_hs__clkbuf_1
X_4775_ _2165_ u_muldiv.o_div\[9\] _2186_ _1913_ VSS VSS VCC VCC _2190_ sky130_fd_sc_hs__a31o_1
X_3726_ u_muldiv.mul\[42\] _1325_ _1452_ VSS VSS VCC VCC _1453_ sky130_fd_sc_hs__a21oi_1
X_3657_ _1106_ csr_data\[5\] _1388_ VSS VSS VCC VCC _1389_ sky130_fd_sc_hs__o21ai_1
X_3588_ _0923_ _1255_ _1272_ VSS VSS VCC VCC _1323_ sky130_fd_sc_hs__a21oi_1
X_5327_ _0917_ _1880_ _2623_ _1841_ VSS VSS VCC VCC _2624_ sky130_fd_sc_hs__a22o_1
X_5258_ _2586_ _2587_ _2590_ _1827_ VSS VSS VCC VCC _2591_ sky130_fd_sc_hs__o211a_1
X_5189_ _2031_ _2105_ _2106_ VSS VSS VCC VCC _2528_ sky130_fd_sc_hs__nor3_1
X_4209_ _1711_ VSS VSS VCC VCC _1778_ sky130_fd_sc_hs__clkbuf_4
X_2890_ _0696_ _0701_ _0704_ VSS VSS VCC VCC _0705_ sky130_fd_sc_hs__o21a_1
X_4560_ _1155_ _2007_ VSS VSS VCC VCC _0273_ sky130_fd_sc_hs__nor2_1
X_4491_ _1976_ VSS VSS VCC VCC _0235_ sky130_fd_sc_hs__clkbuf_1
X_3511_ _0710_ VSS VSS VCC VCC _1248_ sky130_fd_sc_hs__clkinv_2
X_3442_ _1209_ VSS VSS VCC VCC _1210_ sky130_fd_sc_hs__buf_4
X_3373_ _0577_ _1154_ VSS VSS VCC VCC _1155_ sky130_fd_sc_hs__xor2_4
X_5112_ _2039_ _2083_ VSS VSS VCC VCC _2458_ sky130_fd_sc_hs__or2_1
X_5043_ _1305_ _2362_ _2394_ VSS VSS VCC VCC _2395_ sky130_fd_sc_hs__nand3_1
X_4827_ _2181_ _2228_ _2231_ VSS VSS VCC VCC _0316_ sky130_fd_sc_hs__a21oi_1
X_4758_ _2167_ _2176_ u_muldiv.o_div\[5\] VSS VSS VCC VCC _2177_ sky130_fd_sc_hs__a21oi_1
X_4689_ _2109_ _2111_ VSS VSS VCC VCC _2112_ sky130_fd_sc_hs__nand2_1
X_3709_ _0714_ _1435_ _1436_ _0624_ _1145_ VSS VSS VCC VCC _1437_ sky130_fd_sc_hs__o32a_1
Xclkbuf_leaf_32_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_32_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3991_ u_bits.i_op2\[6\] _0688_ _1639_ VSS VSS VCC VCC _1650_ sky130_fd_sc_hs__mux2_1
X_5730_ clknet_leaf_20_i_clk _0373_ VSS VSS VCC VCC u_muldiv.dividend\[14\]
+ sky130_fd_sc_hs__dfxtp_2
X_2942_ u_bits.i_op1\[25\] _0689_ _0649_ VSS VSS VCC VCC _0755_ sky130_fd_sc_hs__mux2_1
X_5661_ clknet_leaf_27_i_clk _0304_ VSS VSS VCC VCC u_muldiv.o_div\[7\] sky130_fd_sc_hs__dfxtp_1
Xclkbuf_leaf_47_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_47_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_2873_ _0687_ VSS VSS VCC VCC _0688_ sky130_fd_sc_hs__buf_4
X_4612_ _2032_ _2033_ _2034_ VSS VSS VCC VCC _2035_ sky130_fd_sc_hs__a21o_1
X_5592_ clknet_leaf_36_i_clk _0239_ VSS VSS VCC VCC u_muldiv.mul\[9\] sky130_fd_sc_hs__dfxtp_1
X_4543_ _2003_ VSS VSS VCC VCC _0260_ sky130_fd_sc_hs__clkbuf_1
X_4474_ _1832_ _1967_ VSS VSS VCC VCC _1968_ sky130_fd_sc_hs__nor2_1
X_3425_ _1192_ _1195_ VSS VSS VCC VCC _1196_ sky130_fd_sc_hs__nand2_1
X_3356_ _1142_ VSS VSS VCC VCC o_add[6] sky130_fd_sc_hs__inv_2
X_3287_ _0644_ _1081_ _0712_ VSS VSS VCC VCC _1082_ sky130_fd_sc_hs__o21a_1
X_5026_ _2379_ VSS VSS VCC VCC _0367_ sky130_fd_sc_hs__clkbuf_1
X_4190_ _1768_ VSS VSS VCC VCC _0142_ sky130_fd_sc_hs__clkbuf_1
X_3210_ _0750_ o_add[27] _0997_ _1010_ _0804_ VSS VSS VCC VCC _1011_ sky130_fd_sc_hs__a221o_1
X_3141_ _0784_ _0780_ _0945_ _0775_ _0825_ _0920_ VSS VSS VCC VCC _0946_ sky130_fd_sc_hs__mux4_2
X_3072_ u_bits.i_op1\[3\] u_bits.i_op1\[2\] _0791_ u_bits.i_op1\[0\] _0657_ _0648_
+ VSS VSS VCC VCC _0881_ sky130_fd_sc_hs__mux4_1
X_3974_ _1595_ VSS VSS VCC VCC _1638_ sky130_fd_sc_hs__clkbuf_4
X_5713_ clknet_leaf_32_i_clk _0356_ VSS VSS VCC VCC u_muldiv.quotient_msk\[27\]
+ sky130_fd_sc_hs__dfxtp_1
X_2925_ _0736_ _0738_ VSS VSS VCC VCC o_add[21] sky130_fd_sc_hs__xnor2_4
X_2856_ _0652_ _0660_ _0664_ _0667_ _0669_ _0670_ VSS VSS VCC VCC _0671_ sky130_fd_sc_hs__mux4_2
X_5644_ clknet_leaf_39_i_clk _0291_ VSS VSS VCC VCC u_muldiv.add_prev\[30\]
+ sky130_fd_sc_hs__dfxtp_1
X_5575_ clknet_leaf_9_i_clk _0222_ VSS VSS VCC VCC u_muldiv.divisor\[56\]
+ sky130_fd_sc_hs__dfxtp_1
X_2787_ _0582_ _0583_ VSS VSS VCC VCC _0602_ sky130_fd_sc_hs__nor2_1
X_4526_ u_muldiv.mul\[22\] u_muldiv.mul\[23\] _1989_ VSS VSS VCC VCC _1995_
+ sky130_fd_sc_hs__mux2_1
X_4457_ u_muldiv.divisor\[57\] _1836_ _1946_ u_muldiv.divisor\[58\] _1954_ VSS VSS
+ VCC VCC _0223_ sky130_fd_sc_hs__a221o_1
X_3408_ _1128_ _1130_ _1137_ _1178_ VSS VSS VCC VCC _1179_ sky130_fd_sc_hs__and4_1
X_4388_ u_bits.i_op2\[12\] _1895_ VSS VSS VCC VCC _1899_ sky130_fd_sc_hs__or2_1
X_3339_ _1125_ _1129_ VSS VSS VCC VCC _1130_ sky130_fd_sc_hs__nand2_4
X_5009_ _1258_ _2362_ _2363_ VSS VSS VCC VCC _2364_ sky130_fd_sc_hs__nand3_1
X_2710_ _0460_ _0524_ u_bits.i_op1\[3\] _0464_ VSS VSS VCC VCC _0525_ sky130_fd_sc_hs__a22o_1
X_3690_ u_bits.i_op2\[8\] _0785_ _1267_ VSS VSS VCC VCC _1419_ sky130_fd_sc_hs__a21oi_1
X_2641_ _0455_ VSS VSS VCC VCC _0456_ sky130_fd_sc_hs__clkbuf_16
X_5360_ clknet_leaf_39_i_clk _0008_ VSS VSS VCC VCC u_muldiv.mul\[56\] sky130_fd_sc_hs__dfxtp_1
X_5291_ u_muldiv.divisor\[6\] _2614_ _2285_ u_muldiv.divisor\[7\] VSS VSS VCC
+ VCC _0397_ sky130_fd_sc_hs__a22o_1
X_4311_ _1207_ VSS VSS VCC VCC _1835_ sky130_fd_sc_hs__buf_4
X_4242_ csr_data\[4\] i_csr_data[4] _1789_ VSS VSS VCC VCC _1795_ sky130_fd_sc_hs__mux2_1
X_4173_ _1759_ VSS VSS VCC VCC _0134_ sky130_fd_sc_hs__clkbuf_1
X_3124_ _0750_ o_add[24] _0907_ _0930_ _0804_ VSS VSS VCC VCC _0931_ sky130_fd_sc_hs__a221o_1
X_3055_ _0860_ _0863_ _0673_ VSS VSS VCC VCC _0864_ sky130_fd_sc_hs__mux2_1
X_3957_ _0702_ i_op1[31] _1621_ VSS VSS VCC VCC _1631_ sky130_fd_sc_hs__mux2_1
X_2908_ _0722_ VSS VSS VCC VCC _0723_ sky130_fd_sc_hs__buf_2
X_3888_ _1593_ VSS VSS VCC VCC _0015_ sky130_fd_sc_hs__clkbuf_1
X_5627_ clknet_leaf_44_i_clk _0274_ VSS VSS VCC VCC u_muldiv.add_prev\[13\]
+ sky130_fd_sc_hs__dfxtp_1
X_2839_ u_bits.i_op1\[15\] VSS VSS VCC VCC _0654_ sky130_fd_sc_hs__buf_4
X_5558_ clknet_leaf_7_i_clk _0205_ VSS VSS VCC VCC u_muldiv.divisor\[39\]
+ sky130_fd_sc_hs__dfxtp_1
X_4509_ u_muldiv.mul\[14\] u_muldiv.mul\[15\] _1978_ VSS VSS VCC VCC _1986_
+ sky130_fd_sc_hs__mux2_1
X_5489_ clknet_leaf_51_i_clk _0137_ VSS VSS VCC VCC o_wdata[7] sky130_fd_sc_hs__dfxtp_4
X_4860_ u_muldiv.o_div\[25\] u_muldiv.o_div\[26\] _2250_ VSS VSS VCC VCC _2258_
+ sky130_fd_sc_hs__or3_1
X_3811_ u_bits.i_op2\[16\] _0653_ _0637_ _1531_ VSS VSS VCC VCC _1532_ sky130_fd_sc_hs__o22a_1
X_4791_ _1835_ _2200_ _2201_ _2202_ VSS VSS VCC VCC _2203_ sky130_fd_sc_hs__a31o_1
X_3742_ _1331_ _1464_ _1466_ _1467_ _1357_ VSS VSS VCC VCC _1468_ sky130_fd_sc_hs__o221a_1
X_3673_ _1402_ _1403_ _1336_ u_pc_sel.i_pc_next\[6\] VSS VSS VCC VCC o_result[6]
+ sky130_fd_sc_hs__a2bb2o_2
X_5412_ clknet_leaf_4_i_clk _0060_ VSS VSS VCC VCC u_bits.i_op2\[3\] sky130_fd_sc_hs__dfxtp_1
X_5343_ _1151_ _2628_ VSS VSS VCC VCC _0435_ sky130_fd_sc_hs__nor2_1
X_5274_ u_muldiv.dividend\[31\] _2601_ _1835_ VSS VSS VCC VCC _2605_ sky130_fd_sc_hs__o21ai_1
X_4225_ _1786_ VSS VSS VCC VCC _0159_ sky130_fd_sc_hs__clkbuf_1
X_4156_ _1750_ VSS VSS VCC VCC _0126_ sky130_fd_sc_hs__clkbuf_1
X_3107_ _0642_ _0625_ _0799_ VSS VSS VCC VCC _0914_ sky130_fd_sc_hs__and3_2
X_4087_ u_pc_sel.i_pc_next\[4\] i_pc_next[4] _1712_ VSS VSS VCC VCC _1716_
+ sky130_fd_sc_hs__mux2_1
X_3038_ _0461_ u_bits.i_op2\[23\] _0465_ u_bits.i_op1\[23\] VSS VSS VCC VCC
+ _0848_ sky130_fd_sc_hs__a22o_1
X_4989_ u_muldiv.dividend\[6\] _2336_ VSS VSS VCC VCC _2345_ sky130_fd_sc_hs__or2_1
X_4010_ _1445_ _1663_ _1651_ i_op2[10] VSS VSS VCC VCC _1664_ sky130_fd_sc_hs__a22o_1
X_4912_ u_muldiv.quotient_msk\[20\] _2282_ _2283_ u_muldiv.quotient_msk\[21\] VSS
+ VSS VCC VCC _0349_ sky130_fd_sc_hs__a22o_1
X_4843_ u_muldiv.o_div\[22\] _2243_ _2244_ VSS VSS VCC VCC _2245_ sky130_fd_sc_hs__mux2_1
X_4774_ _2189_ VSS VSS VCC VCC _0305_ sky130_fd_sc_hs__clkbuf_1
X_3725_ u_muldiv.dividend\[10\] _1326_ _1327_ u_muldiv.o_div\[10\] _1383_ VSS VSS
+ VCC VCC _1452_ sky130_fd_sc_hs__a221o_1
X_3656_ _0731_ VSS VSS VCC VCC _1388_ sky130_fd_sc_hs__clkbuf_2
X_3587_ _1249_ _1317_ _1321_ VSS VSS VCC VCC _1322_ sky130_fd_sc_hs__a21oi_1
X_5326_ _2063_ _2622_ VSS VSS VCC VCC _2623_ sky130_fd_sc_hs__nand2_1
X_5257_ _2288_ _2589_ VSS VSS VCC VCC _2590_ sky130_fd_sc_hs__nand2_1
X_4208_ _1777_ VSS VSS VCC VCC _0151_ sky130_fd_sc_hs__clkbuf_1
X_5188_ _2031_ _2105_ _2106_ _2120_ VSS VSS VCC VCC _2527_ sky130_fd_sc_hs__o22a_1
X_4139_ _1741_ VSS VSS VCC VCC _0118_ sky130_fd_sc_hs__clkbuf_1
X_3510_ _0620_ _1170_ _1246_ _0625_ _0619_ VSS VSS VCC VCC _1247_ sky130_fd_sc_hs__o2111ai_2
X_4490_ u_muldiv.mul\[5\] u_muldiv.mul\[6\] _1584_ VSS VSS VCC VCC _1976_
+ sky130_fd_sc_hs__mux2_1
X_3441_ _1208_ VSS VSS VCC VCC _1209_ sky130_fd_sc_hs__buf_4
X_3372_ _0519_ _1153_ VSS VSS VCC VCC _1154_ sky130_fd_sc_hs__nand2_1
X_5111_ u_muldiv.dividend\[16\] _2444_ VSS VSS VCC VCC _2457_ sky130_fd_sc_hs__xor2_1
X_5042_ u_bits.i_op1\[9\] _2386_ VSS VSS VCC VCC _2394_ sky130_fd_sc_hs__or2_2
X_4826_ _2161_ _2230_ u_muldiv.o_div\[19\] VSS VSS VCC VCC _2231_ sky130_fd_sc_hs__a21oi_1
X_4757_ u_muldiv.quotient_msk\[5\] _2173_ _2156_ VSS VSS VCC VCC _2176_ sky130_fd_sc_hs__mux2_1
X_4688_ _2110_ VSS VSS VCC VCC _2111_ sky130_fd_sc_hs__inv_2
X_3708_ u_bits.i_op2\[9\] _1250_ _1272_ VSS VSS VCC VCC _1436_ sky130_fd_sc_hs__a21oi_1
X_3639_ _0454_ _1368_ _1370_ _1371_ _1357_ VSS VSS VCC VCC _1372_ sky130_fd_sc_hs__o221a_1
X_5309_ u_muldiv.divisor\[21\] _2616_ _2617_ u_muldiv.divisor\[22\] VSS VSS VCC
+ VCC _0412_ sky130_fd_sc_hs__a22o_1
X_3990_ _1641_ _1648_ _1649_ VSS VSS VCC VCC _0061_ sky130_fd_sc_hs__a21o_1
X_2941_ _0752_ _0753_ _0648_ VSS VSS VCC VCC _0754_ sky130_fd_sc_hs__mux2_1
X_5660_ clknet_leaf_27_i_clk _0303_ VSS VSS VCC VCC u_muldiv.o_div\[6\] sky130_fd_sc_hs__dfxtp_1
X_4611_ u_muldiv.dividend\[21\] u_muldiv.divisor\[21\] VSS VSS VCC VCC _2034_
+ sky130_fd_sc_hs__and2b_1
X_2872_ _0642_ VSS VSS VCC VCC _0687_ sky130_fd_sc_hs__buf_2
X_5591_ clknet_leaf_37_i_clk _0238_ VSS VSS VCC VCC u_muldiv.mul\[8\] sky130_fd_sc_hs__dfxtp_1
X_4542_ u_muldiv.mul\[30\] o_add[0] _1583_ VSS VSS VCC VCC _2003_ sky130_fd_sc_hs__mux2_1
X_4473_ u_bits.i_op2\[30\] _1966_ VSS VSS VCC VCC _1967_ sky130_fd_sc_hs__xnor2_1
X_3424_ _1171_ _1194_ VSS VSS VCC VCC _1195_ sky130_fd_sc_hs__xnor2_1
X_3355_ _0561_ _1138_ VSS VSS VCC VCC _1142_ sky130_fd_sc_hs__xor2_4
X_3286_ _0788_ _1080_ _0911_ VSS VSS VCC VCC _1081_ sky130_fd_sc_hs__o21a_1
X_5025_ u_muldiv.dividend\[8\] _2377_ _2378_ VSS VSS VCC VCC _2379_ sky130_fd_sc_hs__mux2_1
X_4809_ u_muldiv.o_div\[15\] _2210_ u_muldiv.o_div\[16\] VSS VSS VCC VCC _2217_
+ sky130_fd_sc_hs__o21ai_1
X_5789_ clknet_leaf_38_i_clk _0431_ VSS VSS VCC VCC u_muldiv.mul\[37\] sky130_fd_sc_hs__dfxtp_1
X_3140_ _0944_ _0870_ _0774_ VSS VSS VCC VCC _0945_ sky130_fd_sc_hs__mux2_1
X_3071_ u_bits.i_op1\[7\] u_bits.i_op1\[6\] u_bits.i_op1\[5\] u_bits.i_op1\[4\] _0657_
+ _0648_ VSS VSS VCC VCC _0880_ sky130_fd_sc_hs__mux4_2
X_5712_ clknet_leaf_32_i_clk _0355_ VSS VSS VCC VCC u_muldiv.quotient_msk\[26\]
+ sky130_fd_sc_hs__dfxtp_1
X_3973_ _1634_ VSS VSS VCC VCC _1637_ sky130_fd_sc_hs__buf_2
X_2924_ _0467_ _0468_ _0737_ VSS VSS VCC VCC _0738_ sky130_fd_sc_hs__a21bo_1
X_2855_ _0524_ VSS VSS VCC VCC _0670_ sky130_fd_sc_hs__buf_4
X_5643_ clknet_leaf_40_i_clk _0290_ VSS VSS VCC VCC u_muldiv.add_prev\[29\]
+ sky130_fd_sc_hs__dfxtp_1
X_5574_ clknet_leaf_9_i_clk _0221_ VSS VSS VCC VCC u_muldiv.divisor\[55\]
+ sky130_fd_sc_hs__dfxtp_1
X_4525_ _1994_ VSS VSS VCC VCC _0251_ sky130_fd_sc_hs__clkbuf_1
X_2786_ _0568_ _0576_ _0600_ VSS VSS VCC VCC _0601_ sky130_fd_sc_hs__a21o_1
X_4456_ _1832_ _1953_ VSS VSS VCC VCC _1954_ sky130_fd_sc_hs__nor2_1
X_3407_ o_add[0] o_add[1] VSS VSS VCC VCC _1178_ sky130_fd_sc_hs__nor2_1
X_4387_ u_muldiv.divisor\[43\] _1867_ _1887_ u_muldiv.divisor\[44\] _1898_ VSS VSS
+ VCC VCC _0209_ sky130_fd_sc_hs__a221o_1
X_3338_ _0532_ _0544_ VSS VSS VCC VCC _1129_ sky130_fd_sc_hs__nand2_1
X_3269_ _1050_ _1065_ _0447_ VSS VSS VCC VCC _1066_ sky130_fd_sc_hs__a21o_1
X_5008_ u_bits.i_op1\[4\] u_bits.i_op1\[5\] u_bits.i_op1\[6\] _2328_ VSS VSS VCC
+ VCC _2363_ sky130_fd_sc_hs__or4_2
Xclkbuf_leaf_31_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_31_i_clk
+ sky130_fd_sc_hs__clkbuf_16
Xclkbuf_leaf_46_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_46_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_2640_ u_muldiv.i_op2_signed alu_ctrl\[2\] VSS VSS VCC VCC _0455_ sky130_fd_sc_hs__nor2_4
X_5290_ _1209_ VSS VSS VCC VCC _2614_ sky130_fd_sc_hs__buf_2
X_4310_ u_muldiv.divisor\[31\] VSS VSS VCC VCC _1834_ sky130_fd_sc_hs__inv_2
X_4241_ _1794_ VSS VSS VCC VCC _0167_ sky130_fd_sc_hs__clkbuf_1
X_4172_ o_wdata[4] i_reg_data2[4] _1756_ VSS VSS VCC VCC _1759_ sky130_fd_sc_hs__mux2_1
X_3123_ _0908_ _0913_ _0929_ _0747_ VSS VSS VCC VCC _0930_ sky130_fd_sc_hs__o31a_1
X_3054_ _0861_ _0862_ _0696_ VSS VSS VCC VCC _0863_ sky130_fd_sc_hs__mux2_1
X_3956_ _1630_ VSS VSS VCC VCC _0046_ sky130_fd_sc_hs__clkbuf_1
X_2907_ _0619_ _0625_ VSS VSS VCC VCC _0722_ sky130_fd_sc_hs__nor2_2
X_3887_ _1214_ _1591_ _1592_ VSS VSS VCC VCC _1593_ sky130_fd_sc_hs__and3_1
X_5626_ clknet_leaf_43_i_clk _0273_ VSS VSS VCC VCC u_muldiv.add_prev\[12\]
+ sky130_fd_sc_hs__dfxtp_1
X_2838_ u_bits.i_op1\[16\] VSS VSS VCC VCC _0653_ sky130_fd_sc_hs__buf_4
X_5557_ clknet_leaf_7_i_clk _0204_ VSS VSS VCC VCC u_muldiv.divisor\[38\]
+ sky130_fd_sc_hs__dfxtp_1
X_2769_ _0582_ _0583_ VSS VSS VCC VCC _0584_ sky130_fd_sc_hs__xor2_4
X_4508_ _1985_ VSS VSS VCC VCC _0243_ sky130_fd_sc_hs__clkbuf_1
X_5488_ clknet_leaf_51_i_clk _0136_ VSS VSS VCC VCC o_wdata[6] sky130_fd_sc_hs__dfxtp_4
X_4439_ u_bits.i_op2\[23\] _1938_ VSS VSS VCC VCC _1940_ sky130_fd_sc_hs__or2_1
X_4790_ u_muldiv.quotient_msk\[12\] u_muldiv.o_div\[12\] _1841_ VSS VSS VCC
+ VCC _2202_ sky130_fd_sc_hs__o21a_1
X_3810_ _0618_ _0639_ _1530_ VSS VSS VCC VCC _1531_ sky130_fd_sc_hs__and3_1
X_3741_ u_muldiv.mul\[11\] _1330_ _1400_ VSS VSS VCC VCC _1467_ sky130_fd_sc_hs__o21ai_1
X_3672_ _1106_ csr_data\[6\] _1388_ VSS VSS VCC VCC _1403_ sky130_fd_sc_hs__o21ai_1
X_5411_ clknet_leaf_49_i_clk _0059_ VSS VSS VCC VCC u_bits.i_op2\[2\] sky130_fd_sc_hs__dfxtp_2
X_5342_ _1145_ _2628_ VSS VSS VCC VCC _0434_ sky130_fd_sc_hs__nor2_1
X_5273_ u_muldiv.dividend\[30\] _2157_ _2604_ VSS VSS VCC VCC _0389_ sky130_fd_sc_hs__a21o_1
X_4224_ u_wr_mux.i_reg_data2\[29\] i_reg_data2[29] _1778_ VSS VSS VCC VCC
+ _1786_ sky130_fd_sc_hs__mux2_1
X_4155_ _0454_ i_alu_ctrl[1] _1745_ VSS VSS VCC VCC _1750_ sky130_fd_sc_hs__mux2_1
X_3106_ _0644_ _0912_ _0712_ VSS VSS VCC VCC _0913_ sky130_fd_sc_hs__o21a_1
X_4086_ _1715_ VSS VSS VCC VCC _0091_ sky130_fd_sc_hs__clkbuf_1
X_3037_ _0739_ csr_data\[22\] _0847_ _0732_ VSS VSS VCC VCC o_result[22] sky130_fd_sc_hs__o211a_2
X_4988_ _2344_ VSS VSS VCC VCC _0364_ sky130_fd_sc_hs__clkbuf_1
X_3939_ _0691_ i_op1[22] _1621_ VSS VSS VCC VCC _1622_ sky130_fd_sc_hs__mux2_1
X_5609_ clknet_leaf_33_i_clk _0256_ VSS VSS VCC VCC u_muldiv.mul\[26\] sky130_fd_sc_hs__dfxtp_1
X_4911_ _1946_ VSS VSS VCC VCC _2283_ sky130_fd_sc_hs__buf_2
X_4842_ _2153_ VSS VSS VCC VCC _2244_ sky130_fd_sc_hs__buf_4
X_4773_ u_muldiv.o_div\[8\] _2188_ _2154_ VSS VSS VCC VCC _2189_ sky130_fd_sc_hs__mux2_1
X_3724_ _0714_ _1449_ _1450_ _0624_ _1151_ VSS VSS VCC VCC _1451_ sky130_fd_sc_hs__o32a_1
X_3655_ _0454_ _1382_ _1385_ _1386_ _1357_ VSS VSS VCC VCC _1387_ sky130_fd_sc_hs__o221a_1
X_3586_ _1265_ _1318_ _1320_ _0906_ VSS VSS VCC VCC _1321_ sky130_fd_sc_hs__o211ai_1
X_5325_ u_muldiv.divisor\[0\] u_muldiv.dividend\[0\] VSS VSS VCC VCC _2622_
+ sky130_fd_sc_hs__or2b_1
X_5256_ _0697_ _2588_ VSS VSS VCC VCC _2589_ sky130_fd_sc_hs__xnor2_1
X_4207_ u_wr_mux.i_reg_data2\[21\] i_reg_data2[21] _1767_ VSS VSS VCC VCC
+ _1777_ sky130_fd_sc_hs__mux2_1
X_5187_ u_muldiv.dividend\[22\] _2506_ u_muldiv.dividend\[23\] VSS VSS VCC VCC
+ _2526_ sky130_fd_sc_hs__o21ai_1
X_4138_ o_pc_target[12] i_pc_target[12] _1734_ VSS VSS VCC VCC _1741_ sky130_fd_sc_hs__mux2_1
X_4069_ u_bits.i_op2\[28\] _1687_ _1596_ i_op2[28] VSS VSS VCC VCC _1705_
+ sky130_fd_sc_hs__a22o_1
X_3440_ _1207_ VSS VSS VCC VCC _1208_ sky130_fd_sc_hs__clkbuf_4
X_3371_ _1152_ _0607_ _0578_ VSS VSS VCC VCC _1153_ sky130_fd_sc_hs__a21o_1
X_5110_ _2456_ VSS VSS VCC VCC _0374_ sky130_fd_sc_hs__clkbuf_1
X_5041_ u_muldiv.dividend\[10\] _2380_ VSS VSS VCC VCC _2393_ sky130_fd_sc_hs__xor2_1
X_4825_ u_muldiv.quotient_msk\[19\] _2226_ _2229_ VSS VSS VCC VCC _2230_ sky130_fd_sc_hs__mux2_1
X_4756_ _2165_ u_muldiv.o_div\[5\] _2173_ _1913_ VSS VSS VCC VCC _2175_ sky130_fd_sc_hs__a31o_1
X_4687_ u_muldiv.divisor\[24\] u_muldiv.dividend\[24\] VSS VSS VCC VCC _2110_
+ sky130_fd_sc_hs__xor2_1
X_3707_ _0908_ _1434_ VSS VSS VCC VCC _1435_ sky130_fd_sc_hs__nor2_1
X_3638_ u_muldiv.mul\[4\] _1330_ _1331_ VSS VSS VCC VCC _1371_ sky130_fd_sc_hs__o21ai_1
X_3569_ _1124_ u_pc_sel.i_pc_next\[1\] _1304_ VSS VSS VCC VCC o_result[1]
+ sky130_fd_sc_hs__o21a_2
X_5308_ u_muldiv.divisor\[20\] _2616_ _2617_ u_muldiv.divisor\[21\] VSS VSS VCC
+ VCC _0411_ sky130_fd_sc_hs__a22o_1
X_5239_ u_muldiv.dividend\[27\] _2164_ _2573_ VSS VSS VCC VCC _0386_ sky130_fd_sc_hs__o21a_1
X_2940_ u_bits.i_op1\[23\] u_bits.i_op1\[24\] _0649_ VSS VSS VCC VCC _0753_
+ sky130_fd_sc_hs__mux2_1
X_2871_ _0634_ _0641_ _0685_ VSS VSS VCC VCC _0686_ sky130_fd_sc_hs__and3_1
X_4610_ u_muldiv.divisor\[20\] u_muldiv.dividend\[20\] VSS VSS VCC VCC _2033_
+ sky130_fd_sc_hs__or2b_1
X_5590_ clknet_leaf_24_i_clk _0237_ VSS VSS VCC VCC u_muldiv.mul\[7\] sky130_fd_sc_hs__dfxtp_1
X_4541_ _2002_ VSS VSS VCC VCC _0259_ sky130_fd_sc_hs__clkbuf_1
X_4472_ u_bits.i_op2\[29\] _1962_ _1845_ VSS VSS VCC VCC _1966_ sky130_fd_sc_hs__o21a_1
X_3423_ _1070_ _1094_ _1101_ _1193_ VSS VSS VCC VCC _1194_ sky130_fd_sc_hs__a31oi_4
X_3354_ _1141_ VSS VSS VCC VCC o_add[7] sky130_fd_sc_hs__inv_2
X_3285_ _0758_ _0823_ _0704_ VSS VSS VCC VCC _1080_ sky130_fd_sc_hs__o21a_1
X_5024_ _2153_ VSS VSS VCC VCC _2378_ sky130_fd_sc_hs__buf_4
X_4808_ _2181_ _2214_ _2216_ VSS VSS VCC VCC _0312_ sky130_fd_sc_hs__a21oi_1
X_5788_ clknet_leaf_38_i_clk _0430_ VSS VSS VCC VCC u_muldiv.mul\[36\] sky130_fd_sc_hs__dfxtp_1
X_4739_ _2153_ VSS VSS VCC VCC _2161_ sky130_fd_sc_hs__clkbuf_4
X_3070_ _0673_ VSS VSS VCC VCC _0879_ sky130_fd_sc_hs__buf_4
X_5711_ clknet_leaf_33_i_clk _0354_ VSS VSS VCC VCC u_muldiv.quotient_msk\[25\]
+ sky130_fd_sc_hs__dfxtp_1
X_3972_ i_inst_branch _1632_ _1636_ u_pc_sel.i_inst_branch VSS VSS VCC VCC
+ _0056_ sky130_fd_sc_hs__a22o_1
X_2923_ _0470_ _0615_ VSS VSS VCC VCC _0737_ sky130_fd_sc_hs__nand2_1
X_2854_ _0668_ VSS VSS VCC VCC _0669_ sky130_fd_sc_hs__clkbuf_4
X_5642_ clknet_leaf_41_i_clk _0289_ VSS VSS VCC VCC u_muldiv.add_prev\[28\]
+ sky130_fd_sc_hs__dfxtp_1
X_5573_ clknet_leaf_9_i_clk _0220_ VSS VSS VCC VCC u_muldiv.divisor\[54\]
+ sky130_fd_sc_hs__dfxtp_1
X_2785_ _0579_ _0599_ VSS VSS VCC VCC _0600_ sky130_fd_sc_hs__or2_1
X_4524_ u_muldiv.mul\[21\] u_muldiv.mul\[22\] _1989_ VSS VSS VCC VCC _1994_
+ sky130_fd_sc_hs__mux2_1
X_4455_ u_bits.i_op2\[26\] _1952_ VSS VSS VCC VCC _1953_ sky130_fd_sc_hs__xnor2_1
X_3406_ _0538_ _0542_ VSS VSS VCC VCC o_add[1] sky130_fd_sc_hs__xor2_4
X_4386_ _1896_ _1897_ VSS VSS VCC VCC _1898_ sky130_fd_sc_hs__nor2_1
X_3337_ _1128_ VSS VSS VCC VCC o_add[3] sky130_fd_sc_hs__inv_2
X_3268_ _0750_ o_add[29] _1063_ _1064_ _0804_ VSS VSS VCC VCC _1065_ sky130_fd_sc_hs__a221o_1
X_5007_ _2293_ VSS VSS VCC VCC _2362_ sky130_fd_sc_hs__buf_2
X_3199_ _0644_ _0999_ _0712_ VSS VSS VCC VCC _1000_ sky130_fd_sc_hs__o21a_1
X_4240_ csr_data\[3\] i_csr_data[3] _1789_ VSS VSS VCC VCC _1794_ sky130_fd_sc_hs__mux2_1
X_4171_ _1758_ VSS VSS VCC VCC _0133_ sky130_fd_sc_hs__clkbuf_1
X_3122_ _0914_ _0921_ _0924_ _0925_ _0928_ VSS VSS VCC VCC _0929_ sky130_fd_sc_hs__a221o_1
X_3053_ _0756_ _0761_ _0663_ VSS VSS VCC VCC _0862_ sky130_fd_sc_hs__mux2_1
X_3955_ _0699_ i_op1[30] _1621_ VSS VSS VCC VCC _1630_ sky130_fd_sc_hs__mux2_1
X_2906_ _0633_ VSS VSS VCC VCC _0721_ sky130_fd_sc_hs__buf_2
X_5625_ clknet_leaf_43_i_clk _0272_ VSS VSS VCC VCC u_muldiv.add_prev\[11\]
+ sky130_fd_sc_hs__dfxtp_1
X_3886_ u_muldiv.i_op2_signed _0626_ _1194_ VSS VSS VCC VCC _1592_ sky130_fd_sc_hs__o21ai_1
X_2837_ _0630_ _0645_ _0646_ _0647_ _0648_ _0651_ VSS VSS VCC VCC _0652_ sky130_fd_sc_hs__mux4_1
X_5556_ clknet_leaf_7_i_clk _0203_ VSS VSS VCC VCC u_muldiv.divisor\[37\]
+ sky130_fd_sc_hs__dfxtp_1
X_2768_ u_bits.i_op1\[11\] u_muldiv.add_prev\[11\] _0450_ VSS VSS VCC VCC
+ _0583_ sky130_fd_sc_hs__mux2_2
X_4507_ u_muldiv.mul\[13\] u_muldiv.mul\[14\] _1978_ VSS VSS VCC VCC _1985_
+ sky130_fd_sc_hs__mux2_1
X_2699_ u_bits.i_op1\[13\] u_muldiv.add_prev\[13\] _0449_ VSS VSS VCC VCC
+ _0514_ sky130_fd_sc_hs__mux2_1
X_5487_ clknet_leaf_51_i_clk _0135_ VSS VSS VCC VCC o_wdata[5] sky130_fd_sc_hs__dfxtp_4
X_4438_ u_bits.i_op2\[23\] _1938_ VSS VSS VCC VCC _1939_ sky130_fd_sc_hs__nand2_1
X_4369_ _1868_ _1883_ u_bits.i_op2\[9\] VSS VSS VCC VCC _1884_ sky130_fd_sc_hs__a21oi_1
X_3740_ u_muldiv.mul\[43\] _1325_ _1465_ VSS VSS VCC VCC _1466_ sky130_fd_sc_hs__a21oi_1
X_3671_ _0454_ _1397_ _1399_ _1401_ _1357_ VSS VSS VCC VCC _1402_ sky130_fd_sc_hs__o221a_1
X_5410_ clknet_leaf_49_i_clk _0058_ VSS VSS VCC VCC u_bits.i_op2\[1\] sky130_fd_sc_hs__dfxtp_1
X_5341_ _1147_ _2628_ VSS VSS VCC VCC _0433_ sky130_fd_sc_hs__nor2_1
X_5272_ _1209_ _2600_ _2603_ _2161_ VSS VSS VCC VCC _2604_ sky130_fd_sc_hs__o211a_1
X_4223_ _1785_ VSS VSS VCC VCC _0158_ sky130_fd_sc_hs__clkbuf_1
X_4154_ _1749_ VSS VSS VCC VCC _0125_ sky130_fd_sc_hs__clkbuf_1
X_3105_ _0909_ _0910_ _0911_ VSS VSS VCC VCC _0912_ sky130_fd_sc_hs__o21a_1
X_4085_ u_pc_sel.i_pc_next\[3\] i_pc_next[3] _1712_ VSS VSS VCC VCC _1715_
+ sky130_fd_sc_hs__mux2_1
X_3036_ _0817_ _0846_ _0447_ VSS VSS VCC VCC _0847_ sky130_fd_sc_hs__a21o_1
Xclkbuf_leaf_30_i_clk clknet_2_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_30_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4987_ u_muldiv.dividend\[5\] _2343_ _2244_ VSS VSS VCC VCC _2344_ sky130_fd_sc_hs__mux2_1
X_3938_ _1595_ VSS VSS VCC VCC _1621_ sky130_fd_sc_hs__clkbuf_4
X_3869_ _1583_ VSS VSS VCC VCC _1584_ sky130_fd_sc_hs__clkbuf_4
Xclkbuf_leaf_45_i_clk clknet_2_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_45_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5608_ clknet_leaf_33_i_clk _0255_ VSS VSS VCC VCC u_muldiv.mul\[25\] sky130_fd_sc_hs__dfxtp_1
X_5539_ clknet_leaf_15_i_clk _0187_ VSS VSS VCC VCC csr_data\[23\] sky130_fd_sc_hs__dfxtp_1
X_4910_ u_muldiv.quotient_msk\[19\] _2282_ _2281_ u_muldiv.quotient_msk\[20\] VSS
+ VSS VCC VCC _0348_ sky130_fd_sc_hs__a22o_1
X_4841_ _2208_ _2240_ _2241_ _2242_ VSS VSS VCC VCC _2243_ sky130_fd_sc_hs__a31o_1
X_4772_ _1835_ _2185_ _2186_ _2187_ VSS VSS VCC VCC _2188_ sky130_fd_sc_hs__a31o_1
X_3723_ _1445_ _1305_ _1272_ VSS VSS VCC VCC _1450_ sky130_fd_sc_hs__a21oi_1
X_3654_ u_muldiv.mul\[5\] _1330_ _1331_ VSS VSS VCC VCC _1386_ sky130_fd_sc_hs__o21ai_1
X_3585_ _0923_ _1255_ _1293_ _1319_ VSS VSS VCC VCC _1320_ sky130_fd_sc_hs__a2bb2o_1
X_5324_ _1913_ _2621_ VSS VSS VCC VCC _0423_ sky130_fd_sc_hs__nor2_1
X_5255_ _0996_ _1029_ _2568_ _2292_ VSS VSS VCC VCC _2588_ sky130_fd_sc_hs__o31a_1
X_4206_ _1776_ VSS VSS VCC VCC _0150_ sky130_fd_sc_hs__clkbuf_1
X_5186_ u_muldiv.dividend\[23\] u_muldiv.dividend\[22\] _2506_ VSS VSS VCC VCC
+ _2525_ sky130_fd_sc_hs__or3_1
X_4137_ _1740_ VSS VSS VCC VCC _0117_ sky130_fd_sc_hs__clkbuf_1
X_4068_ u_bits.i_op2\[29\] u_bits.i_op2\[27\] _1198_ VSS VSS VCC VCC _1704_
+ sky130_fd_sc_hs__mux2_1
X_3019_ _0691_ u_bits.i_op2\[22\] _0637_ _0829_ VSS VSS VCC VCC _0830_ sky130_fd_sc_hs__o22a_1
X_3370_ _0568_ _0576_ _0599_ VSS VSS VCC VCC _1152_ sky130_fd_sc_hs__a21o_1
X_5040_ _2392_ VSS VSS VCC VCC _0368_ sky130_fd_sc_hs__clkbuf_1
X_4824_ _1206_ VSS VSS VCC VCC _2229_ sky130_fd_sc_hs__buf_4
X_4755_ u_muldiv.o_div\[4\] _2171_ _2174_ _2164_ VSS VSS VCC VCC _0301_ sky130_fd_sc_hs__a22o_1
X_3706_ _1110_ _0949_ _1431_ _1249_ _1433_ VSS VSS VCC VCC _1434_ sky130_fd_sc_hs__a221o_1
X_4686_ _2107_ _2108_ VSS VSS VCC VCC _2109_ sky130_fd_sc_hs__nor2_1
X_3637_ u_muldiv.mul\[36\] _1325_ _1369_ VSS VSS VCC VCC _1370_ sky130_fd_sc_hs__a21oi_1
X_3568_ _0446_ csr_data\[1\] _1300_ _1303_ _0730_ VSS VSS VCC VCC _1304_ sky130_fd_sc_hs__a221o_1
X_5307_ u_muldiv.divisor\[19\] _2616_ _2617_ u_muldiv.divisor\[20\] VSS VSS VCC
+ VCC _0410_ sky130_fd_sc_hs__a22o_1
X_3499_ o_wdata[7] _1233_ _0799_ u_wr_mux.i_reg_data2\[15\] VSS VSS VCC VCC
+ _1241_ sky130_fd_sc_hs__a22o_1
X_5238_ _1209_ _2564_ _2565_ _2157_ _2572_ VSS VSS VCC VCC _2573_ sky130_fd_sc_hs__a311o_1
X_5169_ _2508_ _2509_ VSS VSS VCC VCC _2510_ sky130_fd_sc_hs__xnor2_1
X_2870_ _0644_ _0671_ _0684_ VSS VSS VCC VCC _0685_ sky130_fd_sc_hs__o21ai_1
X_4540_ u_muldiv.mul\[29\] u_muldiv.mul\[30\] _1583_ VSS VSS VCC VCC _2002_
+ sky130_fd_sc_hs__mux2_1
X_4471_ u_muldiv.divisor\[60\] _1836_ _1946_ u_muldiv.divisor\[61\] _1965_ VSS VSS
+ VCC VCC _0226_ sky130_fd_sc_hs__a221o_1
X_3422_ _1102_ VSS VSS VCC VCC _1193_ sky130_fd_sc_hs__inv_2
X_3353_ _0556_ _1140_ VSS VSS VCC VCC _1141_ sky130_fd_sc_hs__xnor2_4
X_3284_ u_muldiv.mul\[30\] _0740_ _0720_ u_muldiv.mul\[62\] _1078_ VSS VSS VCC
+ VCC _1079_ sky130_fd_sc_hs__a221o_1
X_5023_ _1878_ _2369_ _2376_ VSS VSS VCC VCC _2377_ sky130_fd_sc_hs__o21a_1
X_4807_ _2167_ _2215_ u_muldiv.o_div\[15\] VSS VSS VCC VCC _2216_ sky130_fd_sc_hs__a21oi_1
X_5787_ clknet_leaf_38_i_clk _0429_ VSS VSS VCC VCC u_muldiv.mul\[35\] sky130_fd_sc_hs__dfxtp_1
X_2999_ _0808_ _0809_ VSS VSS VCC VCC _0811_ sky130_fd_sc_hs__or2_1
X_4738_ _1209_ _2158_ _2159_ _1842_ VSS VSS VCC VCC _2160_ sky130_fd_sc_hs__a31o_1
X_4669_ _2090_ _2091_ VSS VSS VCC VCC _2092_ sky130_fd_sc_hs__and2b_1
X_3971_ i_inst_jal_jalr _1632_ _1636_ u_pc_sel.i_inst_jal_jalr VSS VSS VCC VCC
+ _0055_ sky130_fd_sc_hs__a22o_1
X_5710_ clknet_leaf_33_i_clk _0353_ VSS VSS VCC VCC u_muldiv.quotient_msk\[24\]
+ sky130_fd_sc_hs__dfxtp_1
X_2922_ _0734_ _0735_ VSS VSS VCC VCC _0736_ sky130_fd_sc_hs__xnor2_4
X_2853_ u_bits.i_op2\[2\] VSS VSS VCC VCC _0668_ sky130_fd_sc_hs__clkbuf_4
X_5641_ clknet_leaf_40_i_clk _0288_ VSS VSS VCC VCC u_muldiv.add_prev\[27\]
+ sky130_fd_sc_hs__dfxtp_1
X_2784_ _0590_ _0594_ _0598_ VSS VSS VCC VCC _0599_ sky130_fd_sc_hs__or3_1
X_5572_ clknet_leaf_2_i_clk _0219_ VSS VSS VCC VCC u_muldiv.divisor\[53\]
+ sky130_fd_sc_hs__dfxtp_1
X_4523_ _1993_ VSS VSS VCC VCC _0250_ sky130_fd_sc_hs__clkbuf_1
X_4454_ _1942_ _1951_ _1845_ VSS VSS VCC VCC _1952_ sky130_fd_sc_hs__o21a_1
X_3405_ _0541_ _0540_ VSS VSS VCC VCC o_add[0] sky130_fd_sc_hs__xor2_4
X_4385_ u_bits.i_op2\[12\] _1852_ _1895_ _1856_ VSS VSS VCC VCC _1897_ sky130_fd_sc_hs__a31o_1
X_3336_ _1126_ _1127_ VSS VSS VCC VCC _1128_ sky130_fd_sc_hs__xnor2_4
X_5006_ u_muldiv.dividend\[7\] _2345_ VSS VSS VCC VCC _2361_ sky130_fd_sc_hs__or2_1
X_3267_ _0629_ _1059_ _0955_ VSS VSS VCC VCC _1064_ sky130_fd_sc_hs__a21oi_1
X_3198_ _0909_ _0998_ _0911_ VSS VSS VCC VCC _0999_ sky130_fd_sc_hs__o21a_1
X_4170_ o_wdata[3] i_reg_data2[3] _1756_ VSS VSS VCC VCC _1758_ sky130_fd_sc_hs__mux2_1
X_3121_ _0904_ _0905_ _0926_ _0927_ VSS VSS VCC VCC _0928_ sky130_fd_sc_hs__o22a_1
X_3052_ _0753_ _0755_ _0663_ VSS VSS VCC VCC _0861_ sky130_fd_sc_hs__mux2_1
X_3954_ _1629_ VSS VSS VCC VCC _0045_ sky130_fd_sc_hs__clkbuf_1
X_2905_ _0719_ VSS VSS VCC VCC _0720_ sky130_fd_sc_hs__buf_2
X_3885_ u_muldiv.i_op2_signed _0626_ _1194_ VSS VSS VCC VCC _1591_ sky130_fd_sc_hs__or3_1
X_5624_ clknet_leaf_44_i_clk _0271_ VSS VSS VCC VCC u_muldiv.add_prev\[10\]
+ sky130_fd_sc_hs__dfxtp_1
X_2836_ _0650_ VSS VSS VCC VCC _0651_ sky130_fd_sc_hs__buf_4
X_5555_ clknet_leaf_8_i_clk _0202_ VSS VSS VCC VCC u_muldiv.divisor\[36\]
+ sky130_fd_sc_hs__dfxtp_1
X_2767_ _0456_ _0581_ VSS VSS VCC VCC _0582_ sky130_fd_sc_hs__xnor2_4
X_4506_ _1984_ VSS VSS VCC VCC _0242_ sky130_fd_sc_hs__clkbuf_1
X_2698_ _0456_ _0512_ VSS VSS VCC VCC _0513_ sky130_fd_sc_hs__xnor2_1
X_5486_ clknet_leaf_51_i_clk _0134_ VSS VSS VCC VCC o_wdata[4] sky130_fd_sc_hs__dfxtp_4
X_4437_ u_bits.i_op2\[22\] _1934_ _1846_ VSS VSS VCC VCC _1938_ sky130_fd_sc_hs__o21ai_1
X_4368_ _1406_ u_bits.i_op2\[8\] _1873_ VSS VSS VCC VCC _1883_ sky130_fd_sc_hs__or3_1
X_4299_ _1824_ VSS VSS VCC VCC _0195_ sky130_fd_sc_hs__clkbuf_1
X_3319_ _0783_ VSS VSS VCC VCC _1112_ sky130_fd_sc_hs__buf_4
X_3670_ u_muldiv.mul\[6\] _1330_ _1400_ VSS VSS VCC VCC _1401_ sky130_fd_sc_hs__o21ai_1
X_5340_ _1584_ VSS VSS VCC VCC _2628_ sky130_fd_sc_hs__buf_2
X_5271_ _2601_ _2602_ _1835_ VSS VSS VCC VCC _2603_ sky130_fd_sc_hs__o21ai_1
X_4222_ u_wr_mux.i_reg_data2\[28\] i_reg_data2[28] _1778_ VSS VSS VCC VCC
+ _1785_ sky130_fd_sc_hs__mux2_1
X_4153_ _1639_ i_alu_ctrl[0] _1745_ VSS VSS VCC VCC _1749_ sky130_fd_sc_hs__mux2_1
X_3104_ _0524_ _0703_ VSS VSS VCC VCC _0911_ sky130_fd_sc_hs__nand2_4
X_4084_ _1714_ VSS VSS VCC VCC _0090_ sky130_fd_sc_hs__clkbuf_1
X_3035_ _0750_ o_add[22] _0844_ _0845_ _0804_ VSS VSS VCC VCC _0846_ sky130_fd_sc_hs__a221o_1
X_4986_ _2208_ _2335_ _2336_ _2342_ VSS VSS VCC VCC _2343_ sky130_fd_sc_hs__a31o_1
X_3937_ _1620_ VSS VSS VCC VCC _0037_ sky130_fd_sc_hs__clkbuf_1
X_3868_ _1582_ VSS VSS VCC VCC _1583_ sky130_fd_sc_hs__buf_2
X_3799_ u_muldiv.dividend\[15\] _0742_ _0743_ u_muldiv.o_div\[15\] _0622_ VSS VSS
+ VCC VCC _1521_ sky130_fd_sc_hs__a221o_1
X_5607_ clknet_leaf_33_i_clk _0254_ VSS VSS VCC VCC u_muldiv.mul\[24\] sky130_fd_sc_hs__dfxtp_1
X_2819_ _0620_ _0633_ VSS VSS VCC VCC _0634_ sky130_fd_sc_hs__nand2_2
X_5538_ clknet_leaf_15_i_clk _0186_ VSS VSS VCC VCC csr_data\[22\] sky130_fd_sc_hs__dfxtp_1
X_5469_ clknet_leaf_13_i_clk _0117_ VSS VSS VCC VCC o_pc_target[11] sky130_fd_sc_hs__dfxtp_2
X_4840_ u_muldiv.quotient_msk\[22\] u_muldiv.o_div\[22\] _1840_ VSS VSS VCC
+ VCC _2242_ sky130_fd_sc_hs__o21a_1
X_4771_ u_muldiv.quotient_msk\[8\] u_muldiv.o_div\[8\] _1841_ VSS VSS VCC VCC
+ _2187_ sky130_fd_sc_hs__o21a_1
X_3722_ _0908_ _1448_ VSS VSS VCC VCC _1449_ sky130_fd_sc_hs__nor2_1
X_3653_ u_muldiv.mul\[37\] _1325_ _1384_ VSS VSS VCC VCC _1385_ sky130_fd_sc_hs__a21oi_1
X_5323_ u_muldiv.quotient_msk\[0\] _2152_ u_muldiv.o_div\[0\] VSS VSS VCC VCC
+ _2621_ sky130_fd_sc_hs__a21oi_1
X_3584_ _0923_ _1255_ _0867_ VSS VSS VCC VCC _1319_ sky130_fd_sc_hs__a21o_1
X_5254_ _2030_ _2131_ _2585_ _1839_ VSS VSS VCC VCC _2587_ sky130_fd_sc_hs__a31o_1
X_5185_ _2524_ VSS VSS VCC VCC _0381_ sky130_fd_sc_hs__clkbuf_1
X_4205_ u_wr_mux.i_reg_data2\[20\] i_reg_data2[20] _1767_ VSS VSS VCC VCC
+ _1776_ sky130_fd_sc_hs__mux2_1
X_4136_ o_pc_target[11] i_pc_target[11] _1734_ VSS VSS VCC VCC _1740_ sky130_fd_sc_hs__mux2_1
X_4067_ _1689_ _1702_ _1703_ VSS VSS VCC VCC _0084_ sky130_fd_sc_hs__a21o_1
X_3018_ _0618_ _0639_ _0828_ VSS VSS VCC VCC _0829_ sky130_fd_sc_hs__and3_1
X_4969_ _2068_ _2058_ _2067_ VSS VSS VCC VCC _2327_ sky130_fd_sc_hs__a21o_1
Xclkbuf_leaf_44_i_clk clknet_2_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_44_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4823_ _2170_ u_muldiv.o_div\[19\] _2226_ _2196_ VSS VSS VCC VCC _2228_ sky130_fd_sc_hs__a31o_1
X_4754_ _2165_ _2172_ _2173_ _1842_ u_muldiv.quotient_msk\[4\] VSS VSS VCC VCC
+ _2174_ sky130_fd_sc_hs__a32o_1
X_3705_ u_bits.i_op2\[9\] _1250_ _0926_ _1432_ VSS VSS VCC VCC _1433_ sky130_fd_sc_hs__o22a_1
X_4685_ u_muldiv.dividend\[25\] u_muldiv.divisor\[25\] VSS VSS VCC VCC _2108_
+ sky130_fd_sc_hs__and2b_1
X_3636_ u_muldiv.dividend\[4\] _1326_ _1327_ u_muldiv.o_div\[4\] _0717_ VSS VSS
+ VCC VCC _1369_ sky130_fd_sc_hs__a221o_1
X_3567_ _1301_ _1302_ _0728_ VSS VSS VCC VCC _1303_ sky130_fd_sc_hs__o21a_1
X_5306_ _1842_ VSS VSS VCC VCC _2617_ sky130_fd_sc_hs__buf_2
X_5237_ _2303_ _2567_ _2571_ VSS VSS VCC VCC _2572_ sky130_fd_sc_hs__a21oi_1
X_3498_ _1192_ u_wr_mux.i_reg_data2\[30\] _1240_ VSS VSS VCC VCC o_wdata[30]
+ sky130_fd_sc_hs__a21o_2
X_5168_ _2499_ _2100_ _2033_ VSS VSS VCC VCC _2509_ sky130_fd_sc_hs__o21ai_1
X_5099_ _2444_ _2445_ VSS VSS VCC VCC _2446_ sky130_fd_sc_hs__nand2_1
X_4119_ o_pc_target[3] i_pc_target[3] _1723_ VSS VSS VCC VCC _1731_ sky130_fd_sc_hs__mux2_1
X_4470_ _1963_ _1964_ VSS VSS VCC VCC _1965_ sky130_fd_sc_hs__nor2_1
X_3421_ _0619_ VSS VSS VCC VCC _1192_ sky130_fd_sc_hs__clkbuf_8
X_3352_ _0561_ _1139_ _0570_ VSS VSS VCC VCC _1140_ sky130_fd_sc_hs__o21a_1
X_3283_ u_muldiv.dividend\[30\] _0721_ _0723_ u_muldiv.o_div\[30\] _0744_ VSS VSS
+ VCC VCC _1078_ sky130_fd_sc_hs__a221o_1
X_5022_ _2371_ _2372_ _2374_ _2375_ _1207_ VSS VSS VCC VCC _2376_ sky130_fd_sc_hs__a221o_1
X_4806_ u_muldiv.quotient_msk\[15\] _2210_ _2156_ VSS VSS VCC VCC _2215_ sky130_fd_sc_hs__mux2_1
X_5786_ clknet_leaf_38_i_clk _0428_ VSS VSS VCC VCC u_muldiv.mul\[34\] sky130_fd_sc_hs__dfxtp_1
X_2998_ _0808_ _0809_ VSS VSS VCC VCC _0810_ sky130_fd_sc_hs__nand2_1
X_4737_ u_muldiv.o_div\[2\] _2026_ VSS VSS VCC VCC _2159_ sky130_fd_sc_hs__nand2_1
X_4668_ u_muldiv.divisor\[17\] u_muldiv.dividend\[17\] VSS VSS VCC VCC _2091_
+ sky130_fd_sc_hs__or2b_1
X_3619_ _1274_ _1351_ _1352_ _0624_ _1128_ VSS VSS VCC VCC _1353_ sky130_fd_sc_hs__o32a_1
X_4599_ _1204_ _2023_ VSS VSS VCC VCC _2024_ sky130_fd_sc_hs__nor2_1
X_3970_ i_rd[4] _1632_ _1636_ o_rd[4] VSS VSS VCC VCC _0054_ sky130_fd_sc_hs__a22o_1
X_2921_ u_bits.i_op1\[21\] u_muldiv.add_prev\[21\] _0451_ VSS VSS VCC VCC
+ _0735_ sky130_fd_sc_hs__mux2_2
X_2852_ _0665_ _0666_ _0663_ VSS VSS VCC VCC _0667_ sky130_fd_sc_hs__mux2_1
X_5640_ clknet_leaf_40_i_clk _0287_ VSS VSS VCC VCC u_muldiv.add_prev\[26\]
+ sky130_fd_sc_hs__dfxtp_1
X_2783_ _0596_ _0597_ VSS VSS VCC VCC _0598_ sky130_fd_sc_hs__xnor2_1
X_5571_ clknet_leaf_2_i_clk _0218_ VSS VSS VCC VCC u_muldiv.divisor\[52\]
+ sky130_fd_sc_hs__dfxtp_1
X_4522_ u_muldiv.mul\[20\] u_muldiv.mul\[21\] _1989_ VSS VSS VCC VCC _1993_
+ sky130_fd_sc_hs__mux2_1
X_4453_ _0905_ u_bits.i_op2\[25\] VSS VSS VCC VCC _1951_ sky130_fd_sc_hs__or2_1
X_3404_ o_add[9] o_add[13] o_add[17] VSS VSS VCC VCC _1177_ sky130_fd_sc_hs__or3_1
X_4384_ _1868_ _1895_ u_bits.i_op2\[12\] VSS VSS VCC VCC _1896_ sky130_fd_sc_hs__a21oi_1
X_3335_ _0528_ _0545_ VSS VSS VCC VCC _1127_ sky130_fd_sc_hs__and2b_1
X_3266_ _0628_ _1052_ _1062_ VSS VSS VCC VCC _1063_ sky130_fd_sc_hs__or3_1
X_5005_ u_muldiv.dividend\[7\] _2345_ VSS VSS VCC VCC _2360_ sky130_fd_sc_hs__nand2_1
X_3197_ _0862_ _0859_ _0668_ VSS VSS VCC VCC _0998_ sky130_fd_sc_hs__mux2_1
X_5769_ clknet_leaf_17_i_clk _0412_ VSS VSS VCC VCC u_muldiv.divisor\[21\]
+ sky130_fd_sc_hs__dfxtp_1
X_3120_ _0904_ _0905_ _0867_ VSS VSS VCC VCC _0927_ sky130_fd_sc_hs__a21oi_1
X_3051_ _0704_ _0859_ VSS VSS VCC VCC _0860_ sky130_fd_sc_hs__and2_1
X_3953_ _0697_ i_op1[29] _1621_ VSS VSS VCC VCC _1629_ sky130_fd_sc_hs__mux2_1
X_2904_ _0618_ _0718_ VSS VSS VCC VCC _0719_ sky130_fd_sc_hs__nor2_1
X_3884_ _1590_ VSS VSS VCC VCC _0014_ sky130_fd_sc_hs__clkbuf_1
X_5623_ clknet_leaf_44_i_clk _0270_ VSS VSS VCC VCC u_muldiv.add_prev\[9\]
+ sky130_fd_sc_hs__dfxtp_1
X_2835_ _0649_ VSS VSS VCC VCC _0650_ sky130_fd_sc_hs__buf_4
X_5554_ clknet_leaf_8_i_clk _0201_ VSS VSS VCC VCC u_muldiv.divisor\[35\]
+ sky130_fd_sc_hs__dfxtp_1
X_2766_ _0449_ u_bits.i_op1\[11\] _0497_ _0580_ VSS VSS VCC VCC _0581_ sky130_fd_sc_hs__a31o_1
X_4505_ u_muldiv.mul\[12\] u_muldiv.mul\[13\] _1978_ VSS VSS VCC VCC _1984_
+ sky130_fd_sc_hs__mux2_1
X_2697_ _0449_ u_bits.i_op1\[13\] _0497_ _0511_ VSS VSS VCC VCC _0512_ sky130_fd_sc_hs__a31o_1
X_5485_ clknet_leaf_51_i_clk _0133_ VSS VSS VCC VCC o_wdata[3] sky130_fd_sc_hs__dfxtp_4
X_4436_ u_muldiv.divisor\[53\] _1878_ _1833_ _1936_ _1937_ VSS VSS VCC VCC
+ _0219_ sky130_fd_sc_hs__o221a_1
X_4367_ u_muldiv.divisor\[39\] _1878_ _1829_ u_muldiv.divisor\[40\] _1882_ VSS VSS
+ VCC VCC _0205_ sky130_fd_sc_hs__o221a_1
X_3318_ _0831_ _0699_ _0763_ VSS VSS VCC VCC _1111_ sky130_fd_sc_hs__a21o_1
X_4298_ csr_data\[31\] i_csr_data[31] _1595_ VSS VSS VCC VCC _1824_ sky130_fd_sc_hs__mux2_1
X_3249_ _1045_ _1046_ VSS VSS VCC VCC _1047_ sky130_fd_sc_hs__or2_2
X_5270_ u_muldiv.dividend\[30\] _2583_ VSS VSS VCC VCC _2602_ sky130_fd_sc_hs__and2_1
X_4221_ _1784_ VSS VSS VCC VCC _0157_ sky130_fd_sc_hs__clkbuf_1
X_4152_ _1748_ VSS VSS VCC VCC _0124_ sky130_fd_sc_hs__clkbuf_1
X_3103_ _0690_ _0701_ _0668_ VSS VSS VCC VCC _0910_ sky130_fd_sc_hs__mux2_1
X_4083_ u_pc_sel.i_pc_next\[2\] i_pc_next[2] _1712_ VSS VSS VCC VCC _1714_
+ sky130_fd_sc_hs__mux2_1
X_3034_ _0629_ _0828_ _0714_ VSS VSS VCC VCC _0845_ sky130_fd_sc_hs__a21oi_1
X_4985_ _2229_ _2341_ VSS VSS VCC VCC _2342_ sky130_fd_sc_hs__nor2_1
X_3936_ _0768_ i_op1[21] _1610_ VSS VSS VCC VCC _1620_ sky130_fd_sc_hs__mux2_1
X_3867_ _1198_ u_muldiv.i_on_wait VSS VSS VCC VCC _1582_ sky130_fd_sc_hs__or2_1
X_5606_ clknet_leaf_33_i_clk _0253_ VSS VSS VCC VCC u_muldiv.mul\[23\] sky130_fd_sc_hs__dfxtp_1
X_2818_ _0632_ VSS VSS VCC VCC _0633_ sky130_fd_sc_hs__buf_2
X_3798_ _0714_ _1518_ _1519_ _0623_ _1162_ VSS VSS VCC VCC _1520_ sky130_fd_sc_hs__o32a_1
X_5537_ clknet_leaf_15_i_clk _0185_ VSS VSS VCC VCC csr_data\[21\] sky130_fd_sc_hs__dfxtp_1
X_2749_ _0456_ _0563_ VSS VSS VCC VCC _0564_ sky130_fd_sc_hs__xnor2_4
X_5468_ clknet_leaf_13_i_clk _0116_ VSS VSS VCC VCC o_pc_target[10] sky130_fd_sc_hs__dfxtp_2
X_5399_ clknet_leaf_53_i_clk _0047_ VSS VSS VCC VCC u_bits.i_op1\[31\] sky130_fd_sc_hs__dfxtp_1
X_4419_ u_bits.i_op2\[19\] _1923_ VSS VSS VCC VCC _1924_ sky130_fd_sc_hs__nand2_1
X_4770_ u_muldiv.o_div\[7\] u_muldiv.o_div\[8\] _2179_ VSS VSS VCC VCC _2186_
+ sky130_fd_sc_hs__or3_2
X_3721_ _1110_ _0975_ _1444_ _1248_ _1447_ VSS VSS VCC VCC _1448_ sky130_fd_sc_hs__a221o_1
X_3652_ u_muldiv.dividend\[5\] _1326_ _1327_ u_muldiv.o_div\[5\] _1383_ VSS VSS
+ VCC VCC _1384_ sky130_fd_sc_hs__a221o_1
X_3583_ _0669_ _0788_ _0840_ VSS VSS VCC VCC _1318_ sky130_fd_sc_hs__or3b_1
X_5322_ u_muldiv.outsign _1913_ _2620_ VSS VSS VCC VCC _0422_ sky130_fd_sc_hs__o21a_1
X_5253_ _2030_ _2131_ _2585_ VSS VSS VCC VCC _2586_ sky130_fd_sc_hs__a21oi_1
X_5184_ u_muldiv.dividend\[22\] _2523_ _2485_ VSS VSS VCC VCC _2524_ sky130_fd_sc_hs__mux2_1
X_4204_ _1775_ VSS VSS VCC VCC _0149_ sky130_fd_sc_hs__clkbuf_1
X_4135_ _1739_ VSS VSS VCC VCC _0116_ sky130_fd_sc_hs__clkbuf_1
X_4066_ u_bits.i_op2\[27\] _1687_ _1596_ i_op2[27] VSS VSS VCC VCC _1703_
+ sky130_fd_sc_hs__a22o_1
X_3017_ _0691_ u_bits.i_op2\[22\] VSS VSS VCC VCC _0828_ sky130_fd_sc_hs__nand2_1
X_4968_ _2068_ _2058_ _2067_ VSS VSS VCC VCC _2326_ sky130_fd_sc_hs__nand3_1
X_4899_ _1946_ VSS VSS VCC VCC _2281_ sky130_fd_sc_hs__buf_2
X_3919_ _1611_ VSS VSS VCC VCC _0028_ sky130_fd_sc_hs__clkbuf_1
X_4822_ u_muldiv.o_div\[18\] _2171_ _2227_ _2164_ VSS VSS VCC VCC _0315_ sky130_fd_sc_hs__a22o_1
X_4753_ u_muldiv.o_div\[3\] u_muldiv.o_div\[4\] _2158_ VSS VSS VCC VCC _2173_
+ sky130_fd_sc_hs__or3_2
X_3704_ u_bits.i_op2\[9\] _1250_ _1267_ VSS VSS VCC VCC _1432_ sky130_fd_sc_hs__a21oi_1
X_4684_ u_muldiv.divisor\[25\] u_muldiv.dividend\[25\] VSS VSS VCC VCC _2107_
+ sky130_fd_sc_hs__and2b_1
X_3635_ _1274_ _1366_ _1367_ _0624_ _1137_ VSS VSS VCC VCC _1368_ sky130_fd_sc_hs__o32a_1
X_3566_ u_muldiv.dividend\[1\] _0721_ _0723_ u_muldiv.o_div\[1\] _0724_ VSS VSS
+ VCC VCC _1302_ sky130_fd_sc_hs__a221o_1
X_5305_ u_muldiv.divisor\[18\] _2616_ _2615_ u_muldiv.divisor\[19\] VSS VSS VCC
+ VCC _0409_ sky130_fd_sc_hs__a22o_1
X_3497_ o_wdata[6] _1233_ _0799_ u_wr_mux.i_reg_data2\[14\] VSS VSS VCC VCC
+ _1240_ sky130_fd_sc_hs__a22o_1
X_5236_ _1207_ _2569_ _2570_ _1829_ VSS VSS VCC VCC _2571_ sky130_fd_sc_hs__o31a_1
X_5167_ _2034_ _2032_ VSS VSS VCC VCC _2508_ sky130_fd_sc_hs__and2b_1
X_5098_ u_muldiv.dividend\[14\] _2423_ u_muldiv.dividend\[15\] VSS VSS VCC VCC
+ _2445_ sky130_fd_sc_hs__o21ai_1
X_4118_ _1730_ VSS VSS VCC VCC _0108_ sky130_fd_sc_hs__clkbuf_1
X_4049_ _1689_ _1690_ _1691_ VSS VSS VCC VCC _0078_ sky130_fd_sc_hs__a21o_1
X_3420_ _0618_ _1170_ _1189_ _1190_ _0619_ VSS VSS VCC VCC _1191_ sky130_fd_sc_hs__a221o_1
X_3351_ _1138_ VSS VSS VCC VCC _1139_ sky130_fd_sc_hs__inv_2
X_3282_ _1072_ _1077_ VSS VSS VCC VCC o_add[30] sky130_fd_sc_hs__xor2_4
X_5021_ _1839_ VSS VSS VCC VCC _2375_ sky130_fd_sc_hs__clkbuf_4
X_4805_ _2170_ u_muldiv.o_div\[15\] _2210_ _2196_ VSS VSS VCC VCC _2214_ sky130_fd_sc_hs__a31o_1
X_5785_ clknet_leaf_35_i_clk _0427_ VSS VSS VCC VCC u_muldiv.mul\[33\] sky130_fd_sc_hs__dfxtp_1
X_2997_ u_bits.i_op1\[22\] u_muldiv.add_prev\[22\] _0451_ VSS VSS VCC VCC
+ _0809_ sky130_fd_sc_hs__mux2_1
X_4736_ u_muldiv.o_div\[2\] _2026_ VSS VSS VCC VCC _2158_ sky130_fd_sc_hs__or2_2
X_4667_ u_muldiv.dividend\[17\] u_muldiv.divisor\[17\] VSS VSS VCC VCC _2090_
+ sky130_fd_sc_hs__and2b_1
X_3618_ _0909_ _0794_ _1272_ VSS VSS VCC VCC _1352_ sky130_fd_sc_hs__a21oi_1
X_4598_ op_cnt\[3\] op_cnt\[4\] _2020_ VSS VSS VCC VCC _2023_ sky130_fd_sc_hs__and3_1
X_3549_ _1281_ _1282_ _1283_ _1284_ _0760_ _0879_ VSS VSS VCC VCC _1285_ sky130_fd_sc_hs__mux4_1
X_5219_ u_muldiv.dividend\[25\] _2164_ _2555_ VSS VSS VCC VCC _0384_ sky130_fd_sc_hs__o21ba_1
Xclkbuf_leaf_43_i_clk clknet_2_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_43_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_2920_ _0458_ _0733_ VSS VSS VCC VCC _0734_ sky130_fd_sc_hs__xnor2_4
X_2851_ u_bits.i_op1\[6\] u_bits.i_op1\[5\] _0649_ VSS VSS VCC VCC _0666_
+ sky130_fd_sc_hs__mux2_1
X_2782_ u_bits.i_op1\[8\] u_muldiv.add_prev\[8\] _0450_ VSS VSS VCC VCC _0597_
+ sky130_fd_sc_hs__mux2_1
X_5570_ clknet_leaf_2_i_clk _0217_ VSS VSS VCC VCC u_muldiv.divisor\[51\]
+ sky130_fd_sc_hs__dfxtp_1
X_4521_ _1992_ VSS VSS VCC VCC _0249_ sky130_fd_sc_hs__clkbuf_1
X_4452_ u_muldiv.divisor\[56\] _1836_ _1946_ u_muldiv.divisor\[57\] _1950_ VSS VSS
+ VCC VCC _0222_ sky130_fd_sc_hs__a221o_1
X_3403_ _1176_ VSS VSS VCC VCC o_add[17] sky130_fd_sc_hs__inv_2
X_4383_ _1445_ u_bits.i_op2\[11\] _1888_ VSS VSS VCC VCC _1895_ sky130_fd_sc_hs__or3_1
X_3334_ _0546_ _1125_ VSS VSS VCC VCC _1126_ sky130_fd_sc_hs__nand2_2
X_3265_ _0914_ _1055_ _1058_ _0925_ _1061_ VSS VSS VCC VCC _1062_ sky130_fd_sc_hs__a221o_1
X_5004_ _2356_ _2357_ _2358_ VSS VSS VCC VCC _2359_ sky130_fd_sc_hs__a21oi_1
X_3196_ _0996_ u_bits.i_op2\[27\] _0906_ VSS VSS VCC VCC _0997_ sky130_fd_sc_hs__a21o_1
X_5768_ clknet_leaf_16_i_clk _0411_ VSS VSS VCC VCC u_muldiv.divisor\[20\]
+ sky130_fd_sc_hs__dfxtp_1
X_4719_ u_muldiv.divisor\[55\] u_muldiv.divisor\[54\] u_muldiv.divisor\[53\] u_muldiv.divisor\[52\]
+ VSS VSS VCC VCC _2142_ sky130_fd_sc_hs__or4_1
X_5699_ clknet_leaf_29_i_clk _0342_ VSS VSS VCC VCC u_muldiv.quotient_msk\[13\]
+ sky130_fd_sc_hs__dfxtp_1
X_3050_ u_bits.i_sra _0675_ _0702_ VSS VSS VCC VCC _0859_ sky130_fd_sc_hs__o21a_1
X_3952_ _1628_ VSS VSS VCC VCC _0044_ sky130_fd_sc_hs__clkbuf_1
X_2903_ _0639_ VSS VSS VCC VCC _0718_ sky130_fd_sc_hs__clkbuf_4
X_3883_ o_add[31] _1579_ VSS VSS VCC VCC _1590_ sky130_fd_sc_hs__and2_1
X_5622_ clknet_leaf_44_i_clk _0269_ VSS VSS VCC VCC u_muldiv.add_prev\[8\]
+ sky130_fd_sc_hs__dfxtp_1
X_2834_ u_bits.i_op2\[0\] VSS VSS VCC VCC _0649_ sky130_fd_sc_hs__buf_4
X_5553_ clknet_leaf_8_i_clk _0200_ VSS VSS VCC VCC u_muldiv.divisor\[34\]
+ sky130_fd_sc_hs__dfxtp_1
X_4504_ _1983_ VSS VSS VCC VCC _0241_ sky130_fd_sc_hs__clkbuf_1
X_2765_ _0448_ u_bits.i_op2\[11\] VSS VSS VCC VCC _0580_ sky130_fd_sc_hs__and2b_1
X_2696_ _0448_ u_bits.i_op2\[13\] VSS VSS VCC VCC _0511_ sky130_fd_sc_hs__and2b_1
X_5484_ clknet_leaf_51_i_clk _0132_ VSS VSS VCC VCC o_wdata[2] sky130_fd_sc_hs__dfxtp_4
X_4435_ u_muldiv.divisor\[54\] _1829_ VSS VSS VCC VCC _1937_ sky130_fd_sc_hs__or2_1
X_4366_ u_bits.i_op2\[8\] _1879_ _1881_ VSS VSS VCC VCC _1882_ sky130_fd_sc_hs__a21o_1
X_3317_ _0925_ VSS VSS VCC VCC _1110_ sky130_fd_sc_hs__buf_2
X_4297_ _1823_ VSS VSS VCC VCC _0194_ sky130_fd_sc_hs__clkbuf_1
X_3248_ _1043_ _1044_ VSS VSS VCC VCC _1046_ sky130_fd_sc_hs__nor2_1
X_3179_ _0628_ _0972_ _0981_ VSS VSS VCC VCC _0982_ sky130_fd_sc_hs__or3_2
X_4220_ u_wr_mux.i_reg_data2\[27\] i_reg_data2[27] _1778_ VSS VSS VCC VCC
+ _1784_ sky130_fd_sc_hs__mux2_1
X_4151_ _0618_ i_funct3[2] _1745_ VSS VSS VCC VCC _1748_ sky130_fd_sc_hs__mux2_1
X_3102_ _0788_ VSS VSS VCC VCC _0909_ sky130_fd_sc_hs__buf_4
X_4082_ _1713_ VSS VSS VCC VCC _0089_ sky130_fd_sc_hs__clkbuf_1
X_3033_ _0628_ _0827_ _0830_ _0843_ VSS VSS VCC VCC _0844_ sky130_fd_sc_hs__or4_1
X_4984_ _2337_ _2338_ _2340_ _1826_ VSS VSS VCC VCC _2341_ sky130_fd_sc_hs__o22a_1
X_3935_ _1619_ VSS VSS VCC VCC _0036_ sky130_fd_sc_hs__clkbuf_1
X_5605_ clknet_leaf_33_i_clk _0252_ VSS VSS VCC VCC u_muldiv.mul\[22\] sky130_fd_sc_hs__dfxtp_1
X_3866_ _1581_ VSS VSS VCC VCC _0005_ sky130_fd_sc_hs__clkbuf_1
X_2817_ _0619_ o_funct3[2] VSS VSS VCC VCC _0632_ sky130_fd_sc_hs__and2_1
X_3797_ u_bits.i_op2\[15\] _0654_ _0906_ VSS VSS VCC VCC _1519_ sky130_fd_sc_hs__a21oi_1
X_5536_ clknet_leaf_15_i_clk _0184_ VSS VSS VCC VCC csr_data\[20\] sky130_fd_sc_hs__dfxtp_1
X_2748_ _0459_ u_bits.i_op2\[5\] u_bits.i_op1\[5\] _0463_ VSS VSS VCC VCC
+ _0563_ sky130_fd_sc_hs__a22o_1
X_5467_ clknet_leaf_13_i_clk _0115_ VSS VSS VCC VCC o_pc_target[9] sky130_fd_sc_hs__dfxtp_2
X_2679_ _0488_ _0492_ _0493_ VSS VSS VCC VCC _0494_ sky130_fd_sc_hs__a21o_1
X_4418_ u_bits.i_op2\[18\] _1919_ _1846_ VSS VSS VCC VCC _1923_ sky130_fd_sc_hs__o21ai_1
X_5398_ clknet_leaf_4_i_clk _0046_ VSS VSS VCC VCC u_bits.i_op1\[30\] sky130_fd_sc_hs__dfxtp_2
X_4349_ _1835_ VSS VSS VCC VCC _1867_ sky130_fd_sc_hs__buf_2
X_3720_ _1445_ _1305_ _0926_ _1446_ VSS VSS VCC VCC _1447_ sky130_fd_sc_hs__o22a_1
X_3651_ _0622_ VSS VSS VCC VCC _1383_ sky130_fd_sc_hs__buf_2
X_3582_ _1313_ _1316_ _0644_ VSS VSS VCC VCC _1317_ sky130_fd_sc_hs__mux2_1
X_5321_ _1233_ _1115_ _2618_ _2619_ VSS VSS VCC VCC _2620_ sky130_fd_sc_hs__a31o_1
X_5252_ _2133_ _2132_ VSS VSS VCC VCC _2585_ sky130_fd_sc_hs__and2b_1
X_5183_ _2521_ _2522_ _2229_ VSS VSS VCC VCC _2523_ sky130_fd_sc_hs__mux2_1
X_4203_ u_wr_mux.i_reg_data2\[19\] i_reg_data2[19] _1767_ VSS VSS VCC VCC
+ _1775_ sky130_fd_sc_hs__mux2_1
X_4134_ o_pc_target[10] i_pc_target[10] _1734_ VSS VSS VCC VCC _1739_ sky130_fd_sc_hs__mux2_1
X_4065_ u_bits.i_op2\[28\] u_bits.i_op2\[26\] _1681_ VSS VSS VCC VCC _1702_
+ sky130_fd_sc_hs__mux2_1
X_3016_ _0751_ _0826_ _0712_ VSS VSS VCC VCC _0827_ sky130_fd_sc_hs__o21a_1
X_4967_ _2325_ VSS VSS VCC VCC _0362_ sky130_fd_sc_hs__clkbuf_1
X_4898_ u_muldiv.quotient_msk\[9\] _2280_ _2279_ u_muldiv.quotient_msk\[10\] VSS
+ VSS VCC VCC _0338_ sky130_fd_sc_hs__a22o_1
X_3918_ _0777_ i_op1[12] _1610_ VSS VSS VCC VCC _1611_ sky130_fd_sc_hs__mux2_1
X_3849_ u_muldiv.mul\[19\] _0717_ _0720_ u_muldiv.mul\[51\] _1566_ VSS VSS VCC
+ VCC _1567_ sky130_fd_sc_hs__a221o_1
X_5519_ clknet_leaf_13_i_clk _0167_ VSS VSS VCC VCC csr_data\[3\] sky130_fd_sc_hs__dfxtp_1
X_4821_ _2165_ _2225_ _2226_ _1842_ u_muldiv.quotient_msk\[18\] VSS VSS VCC
+ VCC _2227_ sky130_fd_sc_hs__a32o_1
X_4752_ u_muldiv.o_div\[3\] _2158_ u_muldiv.o_div\[4\] VSS VSS VCC VCC _2172_
+ sky130_fd_sc_hs__o21ai_1
X_4683_ u_muldiv.divisor\[23\] u_muldiv.dividend\[23\] VSS VSS VCC VCC _2106_
+ sky130_fd_sc_hs__and2b_1
X_3703_ _1430_ _1289_ _0940_ _0824_ _0670_ _0643_ VSS VSS VCC VCC _1431_ sky130_fd_sc_hs__mux4_1
X_3634_ _0688_ _1310_ _1272_ VSS VSS VCC VCC _1367_ sky130_fd_sc_hs__a21oi_1
X_3565_ u_muldiv.mul\[1\] _0622_ _0719_ u_muldiv.mul\[33\] VSS VSS VCC VCC
+ _1301_ sky130_fd_sc_hs__a22o_1
X_5304_ u_muldiv.divisor\[17\] _2616_ _2615_ u_muldiv.divisor\[18\] VSS VSS VCC
+ VCC _0408_ sky130_fd_sc_hs__a22o_1
X_3496_ _1192_ u_wr_mux.i_reg_data2\[29\] _1239_ VSS VSS VCC VCC o_wdata[29]
+ sky130_fd_sc_hs__a21o_2
X_5235_ _2362_ _2568_ _0996_ VSS VSS VCC VCC _2570_ sky130_fd_sc_hs__a21oi_1
X_5166_ u_muldiv.dividend\[20\] _2487_ u_muldiv.dividend\[21\] VSS VSS VCC VCC
+ _2507_ sky130_fd_sc_hs__o21ai_1
X_5097_ u_muldiv.dividend\[15\] u_muldiv.dividend\[14\] _2423_ VSS VSS VCC VCC
+ _2444_ sky130_fd_sc_hs__or3_2
X_4117_ o_pc_target[2] i_pc_target[2] _1723_ VSS VSS VCC VCC _1730_ sky130_fd_sc_hs__mux2_1
X_4048_ u_bits.i_op2\[21\] _1687_ _1675_ i_op2[21] VSS VSS VCC VCC _1691_
+ sky130_fd_sc_hs__a22o_1
X_3350_ _1133_ _0566_ _0574_ VSS VSS VCC VCC _1138_ sky130_fd_sc_hs__o21ai_4
X_5020_ _0785_ _2373_ VSS VSS VCC VCC _2374_ sky130_fd_sc_hs__xnor2_1
X_3281_ _1073_ _1075_ _1076_ VSS VSS VCC VCC _1077_ sky130_fd_sc_hs__and3_1
X_4804_ _2213_ VSS VSS VCC VCC _0311_ sky130_fd_sc_hs__clkbuf_1
X_5784_ clknet_leaf_34_i_clk _0426_ VSS VSS VCC VCC u_muldiv.mul\[32\] sky130_fd_sc_hs__dfxtp_1
X_4735_ u_muldiv.outsign _2156_ _2152_ VSS VSS VCC VCC _2157_ sky130_fd_sc_hs__a21oi_4
X_2996_ _0457_ _0807_ VSS VSS VCC VCC _0808_ sky130_fd_sc_hs__xnor2_1
X_4666_ _2087_ _2088_ VSS VSS VCC VCC _2089_ sky130_fd_sc_hs__nand2_1
X_4597_ op_cnt\[3\] _2020_ _2022_ VSS VSS VCC VCC _0295_ sky130_fd_sc_hs__o21a_1
X_3617_ _1249_ _1346_ _1350_ VSS VSS VCC VCC _1351_ sky130_fd_sc_hs__a21oi_1
X_3548_ _1257_ _0786_ u_bits.i_op1\[7\] _0785_ _0778_ _0783_ VSS VSS VCC VCC
+ _1284_ sky130_fd_sc_hs__mux4_1
X_3479_ _1230_ VSS VSS VCC VCC o_wdata[21] sky130_fd_sc_hs__buf_2
X_5218_ _1829_ _2547_ _2554_ _2154_ VSS VSS VCC VCC _2555_ sky130_fd_sc_hs__o211a_1
X_5149_ u_bits.i_op1\[17\] u_bits.i_op1\[18\] _2469_ VSS VSS VCC VCC _2492_
+ sky130_fd_sc_hs__or3_2
X_2850_ u_bits.i_op1\[8\] u_bits.i_op1\[7\] _0649_ VSS VSS VCC VCC _0665_
+ sky130_fd_sc_hs__mux2_1
X_2781_ _0457_ _0595_ VSS VSS VCC VCC _0596_ sky130_fd_sc_hs__xnor2_2
X_4520_ u_muldiv.mul\[20\] u_muldiv.mul\[19\] _1214_ VSS VSS VCC VCC _1992_
+ sky130_fd_sc_hs__mux2_1
X_4451_ _1948_ _1949_ _1833_ VSS VSS VCC VCC _1950_ sky130_fd_sc_hs__a21oi_1
X_3402_ _0610_ _1175_ VSS VSS VCC VCC _1176_ sky130_fd_sc_hs__xor2_2
X_4382_ u_muldiv.divisor\[42\] _1867_ _1887_ u_muldiv.divisor\[43\] _1894_ VSS VSS
+ VCC VCC _0208_ sky130_fd_sc_hs__a221o_1
X_3333_ _0532_ _0544_ VSS VSS VCC VCC _1125_ sky130_fd_sc_hs__or2_1
X_3264_ _0697_ u_bits.i_op2\[29\] _0636_ _1060_ VSS VSS VCC VCC _1061_ sky130_fd_sc_hs__o22a_1
X_5003_ _2356_ _2357_ _1841_ VSS VSS VCC VCC _2358_ sky130_fd_sc_hs__o21ai_1
X_3195_ u_bits.i_op1\[27\] VSS VSS VCC VCC _0996_ sky130_fd_sc_hs__clkbuf_4
X_5767_ clknet_leaf_16_i_clk _0410_ VSS VSS VCC VCC u_muldiv.divisor\[19\]
+ sky130_fd_sc_hs__dfxtp_1
X_2979_ _0791_ u_bits.i_op1\[0\] _0650_ VSS VSS VCC VCC _0792_ sky130_fd_sc_hs__mux2_1
X_5698_ clknet_leaf_29_i_clk _0341_ VSS VSS VCC VCC u_muldiv.quotient_msk\[12\]
+ sky130_fd_sc_hs__dfxtp_1
X_4718_ u_muldiv.divisor\[35\] u_muldiv.divisor\[34\] u_muldiv.divisor\[33\] u_muldiv.divisor\[32\]
+ VSS VSS VCC VCC _2141_ sky130_fd_sc_hs__or4_1
X_4649_ u_muldiv.dividend\[6\] u_muldiv.divisor\[6\] VSS VSS VCC VCC _2072_
+ sky130_fd_sc_hs__and2b_1
X_3951_ _1029_ i_op1[28] _1621_ VSS VSS VCC VCC _1628_ sky130_fd_sc_hs__mux2_1
X_2902_ _0622_ VSS VSS VCC VCC _0717_ sky130_fd_sc_hs__clkbuf_4
X_3882_ _1589_ VSS VSS VCC VCC _0013_ sky130_fd_sc_hs__clkbuf_1
X_5621_ clknet_leaf_46_i_clk _0268_ VSS VSS VCC VCC u_muldiv.add_prev\[7\]
+ sky130_fd_sc_hs__dfxtp_1
X_2833_ _0533_ VSS VSS VCC VCC _0648_ sky130_fd_sc_hs__clkbuf_4
X_5552_ clknet_leaf_8_i_clk _0199_ VSS VSS VCC VCC u_muldiv.divisor\[33\]
+ sky130_fd_sc_hs__dfxtp_1
X_2764_ _0510_ _0577_ _0578_ VSS VSS VCC VCC _0579_ sky130_fd_sc_hs__or3_1
X_4503_ u_muldiv.mul\[11\] u_muldiv.mul\[12\] _1978_ VSS VSS VCC VCC _1983_
+ sky130_fd_sc_hs__mux2_1
X_2695_ _0508_ _0502_ _0509_ VSS VSS VCC VCC _0510_ sky130_fd_sc_hs__or3_1
X_5483_ clknet_leaf_51_i_clk _0131_ VSS VSS VCC VCC o_wdata[1] sky130_fd_sc_hs__dfxtp_4
X_4434_ u_bits.i_op2\[22\] _1935_ VSS VSS VCC VCC _1936_ sky130_fd_sc_hs__xnor2_1
X_4365_ u_bits.i_op2\[8\] _1879_ _1880_ VSS VSS VCC VCC _1881_ sky130_fd_sc_hs__o21ai_1
X_3316_ _0877_ _0882_ _0670_ VSS VSS VCC VCC _1109_ sky130_fd_sc_hs__mux2_1
X_4296_ csr_data\[30\] i_csr_data[30] _1595_ VSS VSS VCC VCC _1823_ sky130_fd_sc_hs__mux2_1
X_3247_ _1043_ _1044_ VSS VSS VCC VCC _1045_ sky130_fd_sc_hs__and2_1
Xclkbuf_leaf_42_i_clk clknet_2_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_42_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3178_ _0914_ _0975_ _0977_ _0925_ _0980_ VSS VSS VCC VCC _0981_ sky130_fd_sc_hs__a221o_1
X_4150_ _1747_ VSS VSS VCC VCC _0123_ sky130_fd_sc_hs__clkbuf_1
X_3101_ _0858_ VSS VSS VCC VCC _0908_ sky130_fd_sc_hs__buf_2
X_4081_ u_pc_sel.i_pc_next\[1\] i_pc_next[1] _1712_ VSS VSS VCC VCC _1713_
+ sky130_fd_sc_hs__mux2_1
X_3032_ _0672_ _0837_ _0842_ _0800_ VSS VSS VCC VCC _0843_ sky130_fd_sc_hs__o211a_1
X_4983_ _1257_ _2339_ VSS VSS VCC VCC _2340_ sky130_fd_sc_hs__xnor2_1
X_3934_ _0630_ i_op1[20] _1610_ VSS VSS VCC VCC _1619_ sky130_fd_sc_hs__mux2_1
X_3865_ o_add[22] _1579_ VSS VSS VCC VCC _1581_ sky130_fd_sc_hs__and2_1
X_5604_ clknet_leaf_33_i_clk _0251_ VSS VSS VCC VCC u_muldiv.mul\[21\] sky130_fd_sc_hs__dfxtp_1
X_2816_ _0630_ u_bits.i_op2\[20\] VSS VSS VCC VCC _0631_ sky130_fd_sc_hs__nand2_1
X_3796_ _1514_ _1517_ VSS VSS VCC VCC _1518_ sky130_fd_sc_hs__nor2_1
X_5535_ clknet_leaf_16_i_clk _0183_ VSS VSS VCC VCC csr_data\[19\] sky130_fd_sc_hs__dfxtp_1
X_2747_ _0556_ _0561_ VSS VSS VCC VCC _0562_ sky130_fd_sc_hs__or2_1
X_5466_ clknet_leaf_13_i_clk _0114_ VSS VSS VCC VCC o_pc_target[8] sky130_fd_sc_hs__dfxtp_2
X_2678_ _0486_ _0487_ VSS VSS VCC VCC _0493_ sky130_fd_sc_hs__nor2_1
X_4417_ u_muldiv.divisor\[49\] _1878_ _1833_ _1921_ _1922_ VSS VSS VCC VCC
+ _0215_ sky130_fd_sc_hs__o221a_1
X_5397_ clknet_leaf_4_i_clk _0045_ VSS VSS VCC VCC u_bits.i_op1\[29\] sky130_fd_sc_hs__dfxtp_1
X_4348_ u_muldiv.divisor\[36\] _1838_ _1843_ u_muldiv.divisor\[37\] _1866_ VSS VSS
+ VCC VCC _0202_ sky130_fd_sc_hs__a221o_1
X_4279_ _1814_ VSS VSS VCC VCC _0185_ sky130_fd_sc_hs__clkbuf_1
X_3650_ _1274_ _1380_ _1381_ _0624_ _1135_ VSS VSS VCC VCC _1382_ sky130_fd_sc_hs__o32a_1
X_3581_ _0970_ _1315_ _0879_ VSS VSS VCC VCC _1316_ sky130_fd_sc_hs__mux2_1
X_5320_ _0619_ _2362_ _1831_ VSS VSS VCC VCC _2619_ sky130_fd_sc_hs__a21o_1
X_5251_ u_muldiv.dividend\[28\] _2564_ u_muldiv.dividend\[29\] VSS VSS VCC VCC
+ _2584_ sky130_fd_sc_hs__o21ai_1
X_4202_ _1774_ VSS VSS VCC VCC _0148_ sky130_fd_sc_hs__clkbuf_1
X_5182_ u_muldiv.dividend\[22\] _2506_ VSS VSS VCC VCC _2522_ sky130_fd_sc_hs__xor2_1
X_4133_ _1738_ VSS VSS VCC VCC _0115_ sky130_fd_sc_hs__clkbuf_1
X_4064_ _1689_ _1700_ _1701_ VSS VSS VCC VCC _0083_ sky130_fd_sc_hs__a21o_1
X_3015_ _0818_ _0822_ _0823_ _0824_ _0825_ _0707_ VSS VSS VCC VCC _0826_ sky130_fd_sc_hs__mux4_2
X_4966_ u_muldiv.dividend\[3\] _2324_ _2244_ VSS VSS VCC VCC _2325_ sky130_fd_sc_hs__mux2_1
X_4897_ u_muldiv.quotient_msk\[8\] _2280_ _2279_ u_muldiv.quotient_msk\[9\] VSS
+ VSS VCC VCC _0337_ sky130_fd_sc_hs__a22o_1
X_3917_ _1595_ VSS VSS VCC VCC _1610_ sky130_fd_sc_hs__clkbuf_4
X_3848_ u_muldiv.dividend\[19\] _0721_ _0723_ u_muldiv.o_div\[19\] _0724_ VSS VSS
+ VCC VCC _1566_ sky130_fd_sc_hs__a221o_1
X_3779_ u_bits.i_op2\[14\] _0655_ _0926_ _1501_ VSS VSS VCC VCC _1502_ sky130_fd_sc_hs__o22a_1
X_5518_ clknet_leaf_13_i_clk _0166_ VSS VSS VCC VCC csr_data\[2\] sky130_fd_sc_hs__dfxtp_1
X_5449_ clknet_leaf_2_i_clk _0097_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[9\]
+ sky130_fd_sc_hs__dfxtp_1
X_4820_ u_muldiv.o_div\[17\] u_muldiv.o_div\[18\] _2218_ VSS VSS VCC VCC _2226_
+ sky130_fd_sc_hs__or3_2
X_4751_ u_muldiv.outsign _2170_ _1913_ VSS VSS VCC VCC _2171_ sky130_fd_sc_hs__a21oi_4
X_4682_ _2035_ _2102_ _2104_ VSS VSS VCC VCC _2105_ sky130_fd_sc_hs__a21oi_1
X_3702_ _1281_ _1282_ _0760_ VSS VSS VCC VCC _1430_ sky130_fd_sc_hs__mux2_1
X_3633_ _1265_ _0681_ _1362_ _1365_ VSS VSS VCC VCC _1366_ sky130_fd_sc_hs__o211a_1
X_3564_ _1298_ _1299_ _0804_ VSS VSS VCC VCC _1300_ sky130_fd_sc_hs__a21o_1
X_5303_ u_muldiv.divisor\[16\] _2616_ _2615_ u_muldiv.divisor\[17\] VSS VSS VCC
+ VCC _0407_ sky130_fd_sc_hs__a22o_1
X_3495_ o_wdata[5] _1233_ _0799_ u_wr_mux.i_reg_data2\[13\] VSS VSS VCC VCC
+ _1239_ sky130_fd_sc_hs__a22o_1
X_5234_ _0996_ _2295_ _2568_ VSS VSS VCC VCC _2569_ sky130_fd_sc_hs__and3_1
X_5165_ u_muldiv.dividend\[21\] u_muldiv.dividend\[20\] _2487_ VSS VSS VCC VCC
+ _2506_ sky130_fd_sc_hs__or3_1
X_4116_ _1729_ VSS VSS VCC VCC _0107_ sky130_fd_sc_hs__clkbuf_1
X_5096_ _2443_ VSS VSS VCC VCC _0373_ sky130_fd_sc_hs__clkbuf_1
X_4047_ u_bits.i_op2\[22\] u_bits.i_op2\[20\] _1681_ VSS VSS VCC VCC _1690_
+ sky130_fd_sc_hs__mux2_1
X_4949_ _1255_ _2293_ _2308_ VSS VSS VCC VCC _2309_ sky130_fd_sc_hs__and3_1
X_3280_ _1021_ _1046_ VSS VSS VCC VCC _1076_ sky130_fd_sc_hs__or2_1
X_4803_ u_muldiv.o_div\[14\] _2212_ _2154_ VSS VSS VCC VCC _2213_ sky130_fd_sc_hs__mux2_1
X_5783_ clknet_leaf_34_i_clk _0425_ VSS VSS VCC VCC u_muldiv.mul\[31\] sky130_fd_sc_hs__dfxtp_1
X_4734_ _1206_ VSS VSS VCC VCC _2156_ sky130_fd_sc_hs__buf_4
X_2995_ _0460_ u_bits.i_op2\[22\] _0464_ u_bits.i_op1\[22\] VSS VSS VCC VCC
+ _0807_ sky130_fd_sc_hs__a22o_1
X_4665_ u_muldiv.dividend\[16\] u_muldiv.divisor\[16\] VSS VSS VCC VCC _2088_
+ sky130_fd_sc_hs__or2b_1
X_4596_ _1204_ _2021_ VSS VSS VCC VCC _2022_ sky130_fd_sc_hs__nor2_1
X_3616_ _1265_ _1347_ _1349_ _0634_ VSS VSS VCC VCC _1350_ sky130_fd_sc_hs__o211ai_1
X_3547_ _0791_ _1255_ _0794_ u_bits.i_op1\[4\] _0651_ _0783_ VSS VSS VCC VCC
+ _1283_ sky130_fd_sc_hs__mux4_1
X_3478_ o_wdata[5] u_wr_mux.i_reg_data2\[21\] _1224_ VSS VSS VCC VCC _1230_
+ sky130_fd_sc_hs__mux2_1
X_5217_ _1831_ _2549_ _2550_ _2553_ _1877_ VSS VSS VCC VCC _2554_ sky130_fd_sc_hs__o32a_1
X_5148_ _2094_ _2489_ _2490_ VSS VSS VCC VCC _2491_ sky130_fd_sc_hs__a21o_1
X_5079_ u_bits.i_op1\[10\] u_bits.i_op1\[11\] u_bits.i_op1\[12\] _2394_ VSS VSS
+ VCC VCC _2428_ sky130_fd_sc_hs__or4_4
X_2780_ _0460_ u_bits.i_op2\[8\] u_bits.i_op1\[8\] _0464_ VSS VSS VCC VCC
+ _0595_ sky130_fd_sc_hs__a22o_1
X_4450_ u_bits.i_op2\[25\] _1947_ VSS VSS VCC VCC _1949_ sky130_fd_sc_hs__or2_1
X_3401_ _0492_ _1164_ VSS VSS VCC VCC _1175_ sky130_fd_sc_hs__nand2_1
X_4381_ _1832_ _1893_ VSS VSS VCC VCC _1894_ sky130_fd_sc_hs__nor2_1
X_3332_ _1106_ csr_data\[31\] _1123_ _1124_ VSS VSS VCC VCC o_result[31] sky130_fd_sc_hs__o211a_2
X_3263_ _0617_ _0638_ _1059_ VSS VSS VCC VCC _1060_ sky130_fd_sc_hs__and3_1
X_5002_ _2073_ _2055_ VSS VSS VCC VCC _2357_ sky130_fd_sc_hs__nor2_1
X_3194_ u_muldiv.mul\[27\] _0740_ _0741_ u_muldiv.mul\[59\] _0994_ VSS VSS VCC
+ VCC _0995_ sky130_fd_sc_hs__a221o_1
X_5766_ clknet_leaf_16_i_clk _0409_ VSS VSS VCC VCC u_muldiv.divisor\[18\]
+ sky130_fd_sc_hs__dfxtp_1
X_2978_ u_bits.i_op1\[1\] VSS VSS VCC VCC _0791_ sky130_fd_sc_hs__clkbuf_4
X_5697_ clknet_leaf_29_i_clk _0340_ VSS VSS VCC VCC u_muldiv.quotient_msk\[11\]
+ sky130_fd_sc_hs__dfxtp_1
X_4717_ u_muldiv.divisor\[43\] u_muldiv.divisor\[42\] u_muldiv.divisor\[41\] _2139_
+ VSS VSS VCC VCC _2140_ sky130_fd_sc_hs__or4_1
X_4648_ _2057_ _2069_ _2070_ VSS VSS VCC VCC _2071_ sky130_fd_sc_hs__o21ba_1
X_4579_ o_add[26] _2004_ VSS VSS VCC VCC _2014_ sky130_fd_sc_hs__and2_1
X_3950_ _1627_ VSS VSS VCC VCC _0043_ sky130_fd_sc_hs__clkbuf_1
X_2901_ _0616_ _0624_ _0715_ VSS VSS VCC VCC _0716_ sky130_fd_sc_hs__o21ai_1
X_3881_ o_add[30] _1579_ VSS VSS VCC VCC _1589_ sky130_fd_sc_hs__and2_1
X_5620_ clknet_leaf_46_i_clk _0267_ VSS VSS VCC VCC u_muldiv.add_prev\[6\]
+ sky130_fd_sc_hs__dfxtp_1
X_2832_ u_bits.i_op1\[17\] VSS VSS VCC VCC _0647_ sky130_fd_sc_hs__buf_4
X_5551_ clknet_leaf_8_i_clk _0198_ VSS VSS VCC VCC u_muldiv.divisor\[32\]
+ sky130_fd_sc_hs__dfxtp_1
X_2763_ _0517_ _0518_ VSS VSS VCC VCC _0578_ sky130_fd_sc_hs__xnor2_1
X_4502_ _1982_ VSS VSS VCC VCC _0240_ sky130_fd_sc_hs__clkbuf_1
X_5482_ clknet_leaf_51_i_clk _0130_ VSS VSS VCC VCC o_wdata[0] sky130_fd_sc_hs__dfxtp_4
X_2694_ _0505_ _0506_ VSS VSS VCC VCC _0509_ sky130_fd_sc_hs__xnor2_4
X_4433_ _1850_ _1934_ VSS VSS VCC VCC _1935_ sky130_fd_sc_hs__nand2_1
X_4364_ u_muldiv.on_wait u_muldiv.i_on_end VSS VSS VCC VCC _1880_ sky130_fd_sc_hs__nor2_4
X_4295_ _1822_ VSS VSS VCC VCC _0193_ sky130_fd_sc_hs__clkbuf_1
X_3315_ u_muldiv.mul\[31\] _0740_ _0720_ u_muldiv.mul\[63\] _1107_ VSS VSS VCC
+ VCC _1108_ sky130_fd_sc_hs__a221o_1
X_3246_ _0697_ u_muldiv.add_prev\[29\] _0452_ VSS VSS VCC VCC _1044_ sky130_fd_sc_hs__mux2_1
X_3177_ _0689_ u_bits.i_op2\[26\] _0636_ _0979_ VSS VSS VCC VCC _0980_ sky130_fd_sc_hs__o22a_1
X_5749_ clknet_leaf_24_i_clk _0392_ VSS VSS VCC VCC u_muldiv.divisor\[1\]
+ sky130_fd_sc_hs__dfxtp_1
X_3100_ _0904_ _0905_ _0906_ VSS VSS VCC VCC _0907_ sky130_fd_sc_hs__a21o_1
X_4080_ _1711_ VSS VSS VCC VCC _1712_ sky130_fd_sc_hs__clkbuf_4
X_3031_ _0674_ _0841_ _0642_ VSS VSS VCC VCC _0842_ sky130_fd_sc_hs__a21bo_1
X_4982_ _1310_ _2328_ _2292_ VSS VSS VCC VCC _2339_ sky130_fd_sc_hs__o21a_1
X_3933_ _1618_ VSS VSS VCC VCC _0035_ sky130_fd_sc_hs__clkbuf_1
X_3864_ _1580_ VSS VSS VCC VCC _0004_ sky130_fd_sc_hs__clkbuf_1
X_5603_ clknet_leaf_33_i_clk _0250_ VSS VSS VCC VCC u_muldiv.mul\[20\] sky130_fd_sc_hs__dfxtp_1
X_2815_ u_bits.i_op1\[20\] VSS VSS VCC VCC _0630_ sky130_fd_sc_hs__buf_4
X_3795_ _1110_ _1109_ _1516_ _0858_ VSS VSS VCC VCC _1517_ sky130_fd_sc_hs__a211o_1
X_5534_ clknet_leaf_14_i_clk _0182_ VSS VSS VCC VCC csr_data\[18\] sky130_fd_sc_hs__dfxtp_1
X_2746_ _0559_ _0560_ VSS VSS VCC VCC _0561_ sky130_fd_sc_hs__xnor2_4
X_5465_ clknet_leaf_13_i_clk _0113_ VSS VSS VCC VCC o_pc_target[7] sky130_fd_sc_hs__dfxtp_2
X_2677_ _0490_ _0491_ VSS VSS VCC VCC _0492_ sky130_fd_sc_hs__nand2_1
X_4416_ u_muldiv.divisor\[50\] _1829_ VSS VSS VCC VCC _1922_ sky130_fd_sc_hs__or2_1
X_5396_ clknet_leaf_4_i_clk _0044_ VSS VSS VCC VCC u_bits.i_op1\[28\] sky130_fd_sc_hs__dfxtp_2
X_4347_ _1864_ _1865_ _1833_ VSS VSS VCC VCC _1866_ sky130_fd_sc_hs__a21oi_1
X_4278_ csr_data\[21\] i_csr_data[21] _1811_ VSS VSS VCC VCC _1814_ sky130_fd_sc_hs__mux2_1
X_3229_ _0687_ _1027_ _0711_ VSS VSS VCC VCC _1028_ sky130_fd_sc_hs__o21a_1
X_3580_ _1314_ _0818_ _0758_ VSS VSS VCC VCC _1315_ sky130_fd_sc_hs__mux2_1
Xclkbuf_leaf_41_i_clk clknet_2_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_41_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5250_ u_muldiv.dividend\[29\] u_muldiv.dividend\[28\] _2564_ VSS VSS VCC VCC
+ _2583_ sky130_fd_sc_hs__or3_1
X_4201_ u_wr_mux.i_reg_data2\[18\] i_reg_data2[18] _1767_ VSS VSS VCC VCC
+ _1774_ sky130_fd_sc_hs__mux2_1
X_5181_ _2105_ _2518_ _2520_ _2375_ VSS VSS VCC VCC _2521_ sky130_fd_sc_hs__a2bb2o_1
X_4132_ o_pc_target[9] i_pc_target[9] _1734_ VSS VSS VCC VCC _1738_ sky130_fd_sc_hs__mux2_1
X_4063_ u_bits.i_op2\[26\] _1687_ _1596_ i_op2[26] VSS VSS VCC VCC _1701_
+ sky130_fd_sc_hs__a22o_1
X_3014_ _0696_ VSS VSS VCC VCC _0825_ sky130_fd_sc_hs__buf_4
X_4965_ _2208_ _2315_ _2316_ _2323_ VSS VSS VCC VCC _2324_ sky130_fd_sc_hs__a31o_1
X_3916_ _1609_ VSS VSS VCC VCC _0027_ sky130_fd_sc_hs__clkbuf_1
X_4896_ u_muldiv.quotient_msk\[7\] _2280_ _2279_ u_muldiv.quotient_msk\[8\] VSS
+ VSS VCC VCC _0336_ sky130_fd_sc_hs__a22o_1
X_3847_ _1106_ csr_data\[18\] _1565_ _1124_ VSS VSS VCC VCC o_result[18] sky130_fd_sc_hs__o211a_2
X_3778_ u_bits.i_op2\[14\] _0655_ _1267_ VSS VSS VCC VCC _1501_ sky130_fd_sc_hs__a21oi_1
X_5517_ clknet_leaf_13_i_clk _0165_ VSS VSS VCC VCC csr_data\[1\] sky130_fd_sc_hs__dfxtp_1
X_2729_ _0538_ _0542_ _0543_ VSS VSS VCC VCC _0544_ sky130_fd_sc_hs__a21oi_1
X_5448_ clknet_leaf_9_i_clk _0096_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[8\]
+ sky130_fd_sc_hs__dfxtp_1
X_5379_ clknet_leaf_47_i_clk _0027_ VSS VSS VCC VCC u_bits.i_op1\[11\] sky130_fd_sc_hs__dfxtp_2
Xclkbuf_2_0__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_0__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4750_ _2156_ VSS VSS VCC VCC _2170_ sky130_fd_sc_hs__clkbuf_4
X_4681_ _2031_ _2103_ VSS VSS VCC VCC _2104_ sky130_fd_sc_hs__or2_1
X_3701_ _1428_ _1429_ _1336_ u_pc_sel.i_pc_next\[8\] VSS VSS VCC VCC o_result[8]
+ sky130_fd_sc_hs__a2bb2o_2
X_3632_ _0858_ _1364_ VSS VSS VCC VCC _1365_ sky130_fd_sc_hs__nor2_1
X_5302_ _1209_ VSS VSS VCC VCC _2616_ sky130_fd_sc_hs__buf_2
X_3563_ _1112_ _0791_ _0906_ _0955_ VSS VSS VCC VCC _1299_ sky130_fd_sc_hs__a211o_1
X_3494_ _1192_ u_wr_mux.i_reg_data2\[28\] _1238_ VSS VSS VCC VCC o_wdata[28]
+ sky130_fd_sc_hs__a21o_2
X_5233_ _0943_ _0689_ _2548_ VSS VSS VCC VCC _2568_ sky130_fd_sc_hs__or3_1
X_5164_ _2505_ VSS VSS VCC VCC _0379_ sky130_fd_sc_hs__clkbuf_1
X_4115_ o_pc_target[1] i_pc_target[1] _1723_ VSS VSS VCC VCC _1729_ sky130_fd_sc_hs__mux2_1
X_5095_ u_muldiv.dividend\[14\] _2442_ _2378_ VSS VSS VCC VCC _2443_ sky130_fd_sc_hs__mux2_1
X_4046_ _1635_ VSS VSS VCC VCC _1689_ sky130_fd_sc_hs__buf_2
X_4948_ u_bits.i_op1\[0\] u_bits.i_op1\[1\] VSS VSS VCC VCC _2308_ sky130_fd_sc_hs__or2_2
X_4879_ u_muldiv.quotient_msk\[30\] u_muldiv.o_div\[30\] VSS VSS VCC VCC _2273_
+ sky130_fd_sc_hs__or2_1
X_4802_ _2208_ _2209_ _2210_ _2211_ VSS VSS VCC VCC _2212_ sky130_fd_sc_hs__a31o_1
X_5782_ clknet_leaf_24_i_clk _0424_ VSS VSS VCC VCC u_muldiv.dividend\[0\]
+ sky130_fd_sc_hs__dfxtp_1
X_2994_ _0739_ csr_data\[21\] _0806_ _0732_ VSS VSS VCC VCC o_result[21] sky130_fd_sc_hs__o211a_2
X_4733_ _2155_ VSS VSS VCC VCC _0298_ sky130_fd_sc_hs__clkbuf_1
X_4664_ u_muldiv.divisor\[16\] u_muldiv.dividend\[16\] VSS VSS VCC VCC _2087_
+ sky130_fd_sc_hs__or2b_1
X_4595_ op_cnt\[3\] _2020_ VSS VSS VCC VCC _2021_ sky130_fd_sc_hs__and2_1
X_3615_ _0909_ _0794_ _1293_ _1348_ VSS VSS VCC VCC _1349_ sky130_fd_sc_hs__a2bb2o_1
X_3546_ u_bits.i_op1\[13\] _0655_ _0654_ _0653_ _0658_ _0779_ VSS VSS VCC VCC
+ _1282_ sky130_fd_sc_hs__mux4_2
X_5216_ _2551_ _2552_ VSS VSS VCC VCC _2553_ sky130_fd_sc_hs__nand2_1
X_3477_ _1229_ VSS VSS VCC VCC o_wdata[20] sky130_fd_sc_hs__buf_2
X_5147_ _2094_ _2489_ _1826_ VSS VSS VCC VCC _2490_ sky130_fd_sc_hs__o21ai_1
X_5078_ _2044_ _2415_ _2425_ _2288_ VSS VSS VCC VCC _2427_ sky130_fd_sc_hs__a31o_1
X_4029_ u_bits.i_op2\[17\] u_bits.i_op2\[15\] _1657_ VSS VSS VCC VCC _1677_
+ sky130_fd_sc_hs__mux2_1
X_3400_ _0612_ _1174_ VSS VSS VCC VCC o_add[16] sky130_fd_sc_hs__xnor2_4
X_4380_ u_bits.i_op2\[11\] _1892_ VSS VSS VCC VCC _1893_ sky130_fd_sc_hs__xnor2_1
X_3331_ _0731_ VSS VSS VCC VCC _1124_ sky130_fd_sc_hs__buf_2
X_3262_ _0697_ u_bits.i_op2\[29\] VSS VSS VCC VCC _1059_ sky130_fd_sc_hs__nand2_1
X_5001_ _2056_ _2348_ VSS VSS VCC VCC _2356_ sky130_fd_sc_hs__or2b_1
X_3193_ u_muldiv.dividend\[27\] _0742_ _0743_ u_muldiv.o_div\[27\] _0744_ VSS VSS
+ VCC VCC _0994_ sky130_fd_sc_hs__a221o_1
X_5765_ clknet_leaf_18_i_clk _0408_ VSS VSS VCC VCC u_muldiv.divisor\[17\]
+ sky130_fd_sc_hs__dfxtp_1
X_2977_ _0775_ _0780_ _0784_ _0787_ _0788_ _0789_ VSS VSS VCC VCC _0790_ sky130_fd_sc_hs__mux4_1
X_5696_ clknet_leaf_29_i_clk _0339_ VSS VSS VCC VCC u_muldiv.quotient_msk\[10\]
+ sky130_fd_sc_hs__dfxtp_1
X_4716_ u_muldiv.divisor\[39\] u_muldiv.divisor\[38\] u_muldiv.divisor\[37\] u_muldiv.divisor\[36\]
+ VSS VSS VCC VCC _2139_ sky130_fd_sc_hs__or4_1
X_4647_ u_muldiv.divisor\[5\] u_muldiv.dividend\[5\] VSS VSS VCC VCC _2070_
+ sky130_fd_sc_hs__and2b_1
X_4578_ _2013_ VSS VSS VCC VCC _0285_ sky130_fd_sc_hs__clkbuf_1
X_3529_ _0916_ _0788_ _0917_ VSS VSS VCC VCC _1266_ sky130_fd_sc_hs__or3b_1
X_2900_ _0629_ _0631_ _0686_ _0713_ _0714_ VSS VSS VCC VCC _0715_ sky130_fd_sc_hs__a221o_1
X_3880_ _1588_ VSS VSS VCC VCC _0012_ sky130_fd_sc_hs__clkbuf_1
X_2831_ u_bits.i_op1\[19\] VSS VSS VCC VCC _0646_ sky130_fd_sc_hs__buf_4
X_5550_ clknet_leaf_8_i_clk _0197_ VSS VSS VCC VCC u_muldiv.divisor\[31\]
+ sky130_fd_sc_hs__dfxtp_1
X_2762_ _0515_ _0520_ VSS VSS VCC VCC _0577_ sky130_fd_sc_hs__or2b_2
X_4501_ u_muldiv.mul\[10\] u_muldiv.mul\[11\] _1978_ VSS VSS VCC VCC _1982_
+ sky130_fd_sc_hs__mux2_1
X_5481_ clknet_leaf_38_i_clk _0129_ VSS VSS VCC VCC u_mux.i_add_override sky130_fd_sc_hs__dfxtp_1
X_2693_ _0500_ _0501_ VSS VSS VCC VCC _0508_ sky130_fd_sc_hs__and2_1
X_4432_ u_bits.i_op2\[21\] u_bits.i_op2\[20\] _1927_ VSS VSS VCC VCC _1934_
+ sky130_fd_sc_hs__or3_1
X_4363_ _1406_ _1873_ _1846_ VSS VSS VCC VCC _1879_ sky130_fd_sc_hs__o21ai_1
X_3314_ u_muldiv.dividend\[31\] _0721_ _0723_ u_muldiv.o_div\[31\] _0724_ VSS VSS
+ VCC VCC _1107_ sky130_fd_sc_hs__a221o_1
X_4294_ csr_data\[29\] i_csr_data[29] _1595_ VSS VSS VCC VCC _1822_ sky130_fd_sc_hs__mux2_1
X_3245_ _0458_ _1042_ VSS VSS VCC VCC _1043_ sky130_fd_sc_hs__xnor2_1
X_3176_ _0617_ _0638_ _0978_ VSS VSS VCC VCC _0979_ sky130_fd_sc_hs__and3_1
X_5748_ clknet_leaf_24_i_clk _0391_ VSS VSS VCC VCC u_muldiv.divisor\[0\]
+ sky130_fd_sc_hs__dfxtp_1
X_5679_ clknet_leaf_31_i_clk _0322_ VSS VSS VCC VCC u_muldiv.o_div\[25\] sky130_fd_sc_hs__dfxtp_1
X_3030_ _0838_ _0840_ _0760_ VSS VSS VCC VCC _0841_ sky130_fd_sc_hs__mux2_1
X_4981_ _2070_ _2057_ _2069_ _1826_ VSS VSS VCC VCC _2338_ sky130_fd_sc_hs__o31ai_1
X_3932_ _0646_ i_op1[19] _1610_ VSS VSS VCC VCC _1618_ sky130_fd_sc_hs__mux2_1
X_3863_ o_add[21] _1579_ VSS VSS VCC VCC _1580_ sky130_fd_sc_hs__and2_1
X_5602_ clknet_leaf_32_i_clk _0249_ VSS VSS VCC VCC u_muldiv.mul\[19\] sky130_fd_sc_hs__dfxtp_1
X_2814_ _0628_ VSS VSS VCC VCC _0629_ sky130_fd_sc_hs__buf_2
X_5533_ clknet_leaf_14_i_clk _0181_ VSS VSS VCC VCC csr_data\[17\] sky130_fd_sc_hs__dfxtp_1
X_3794_ u_bits.i_op2\[15\] _0654_ _0637_ _1515_ VSS VSS VCC VCC _1516_ sky130_fd_sc_hs__o22a_1
X_2745_ u_bits.i_op1\[6\] u_muldiv.add_prev\[6\] _0448_ VSS VSS VCC VCC _0560_
+ sky130_fd_sc_hs__mux2_2
X_5464_ clknet_leaf_14_i_clk _0112_ VSS VSS VCC VCC o_pc_target[6] sky130_fd_sc_hs__dfxtp_2
X_2676_ u_bits.i_op1\[16\] u_muldiv.add_prev\[16\] _0451_ VSS VSS VCC VCC
+ _0491_ sky130_fd_sc_hs__mux2_1
X_5395_ clknet_leaf_53_i_clk _0043_ VSS VSS VCC VCC u_bits.i_op1\[27\] sky130_fd_sc_hs__dfxtp_4
X_4415_ u_bits.i_op2\[18\] _1920_ VSS VSS VCC VCC _1921_ sky130_fd_sc_hs__xnor2_1
X_4346_ _1376_ _1863_ VSS VSS VCC VCC _1865_ sky130_fd_sc_hs__or2_1
X_4277_ _1813_ VSS VSS VCC VCC _0184_ sky130_fd_sc_hs__clkbuf_1
X_3228_ _0788_ _0705_ _0911_ VSS VSS VCC VCC _1027_ sky130_fd_sc_hs__o21a_1
X_3159_ _0960_ _0961_ VSS VSS VCC VCC _0963_ sky130_fd_sc_hs__or2_1
X_4200_ _1773_ VSS VSS VCC VCC _0147_ sky130_fd_sc_hs__clkbuf_1
X_5180_ _0691_ _2519_ VSS VSS VCC VCC _2520_ sky130_fd_sc_hs__xnor2_1
X_4131_ _1737_ VSS VSS VCC VCC _0114_ sky130_fd_sc_hs__clkbuf_1
X_4062_ u_bits.i_op2\[27\] u_bits.i_op2\[25\] _1681_ VSS VSS VCC VCC _1700_
+ sky130_fd_sc_hs__mux2_1
X_3013_ _0703_ VSS VSS VCC VCC _0824_ sky130_fd_sc_hs__inv_2
X_4964_ _2319_ _2320_ _2322_ _2303_ _1827_ VSS VSS VCC VCC _2323_ sky130_fd_sc_hs__o221a_1
X_3915_ _1251_ i_op1[11] _1599_ VSS VSS VCC VCC _1609_ sky130_fd_sc_hs__mux2_1
X_4895_ _1209_ VSS VSS VCC VCC _2280_ sky130_fd_sc_hs__buf_2
X_3846_ _1554_ _1564_ _0446_ VSS VSS VCC VCC _1565_ sky130_fd_sc_hs__a21o_1
X_3777_ _1499_ _1081_ _0643_ VSS VSS VCC VCC _1500_ sky130_fd_sc_hs__mux2_1
X_5516_ clknet_leaf_13_i_clk _0164_ VSS VSS VCC VCC csr_data\[0\] sky130_fd_sc_hs__dfxtp_1
X_2728_ _0536_ _0537_ VSS VSS VCC VCC _0543_ sky130_fd_sc_hs__and2_1
X_5447_ clknet_leaf_2_i_clk _0095_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[7\]
+ sky130_fd_sc_hs__dfxtp_1
X_2659_ _0472_ _0473_ VSS VSS VCC VCC _0474_ sky130_fd_sc_hs__nor2_1
X_5378_ clknet_leaf_47_i_clk _0026_ VSS VSS VCC VCC u_bits.i_op1\[10\] sky130_fd_sc_hs__dfxtp_2
X_4329_ _0915_ _1850_ _0923_ VSS VSS VCC VCC _1851_ sky130_fd_sc_hs__a21oi_1
X_3700_ _1333_ csr_data\[8\] _1388_ VSS VSS VCC VCC _1429_ sky130_fd_sc_hs__o21ai_1
X_4680_ u_muldiv.dividend\[22\] u_muldiv.divisor\[22\] VSS VSS VCC VCC _2103_
+ sky130_fd_sc_hs__and2b_1
X_3631_ _0672_ _1310_ _0637_ _1363_ VSS VSS VCC VCC _1364_ sky130_fd_sc_hs__o22a_1
X_3562_ _0749_ o_add[1] _1297_ _0747_ VSS VSS VCC VCC _1298_ sky130_fd_sc_hs__a22o_1
X_5301_ u_muldiv.divisor\[15\] _2614_ _2615_ u_muldiv.divisor\[16\] VSS VSS VCC
+ VCC _0406_ sky130_fd_sc_hs__a22o_1
X_3493_ o_wdata[4] _1233_ _0799_ u_wr_mux.i_reg_data2\[12\] VSS VSS VCC VCC
+ _1238_ sky130_fd_sc_hs__a22o_1
X_5232_ _2113_ _2566_ VSS VSS VCC VCC _2567_ sky130_fd_sc_hs__xor2_1
X_5163_ u_muldiv.dividend\[20\] _2504_ _2485_ VSS VSS VCC VCC _2505_ sky130_fd_sc_hs__mux2_1
X_4114_ i_res_src[2] _1638_ _1635_ o_res_src[2] VSS VSS VCC VCC _0106_ sky130_fd_sc_hs__a22o_1
X_5094_ _2435_ _2441_ _1877_ VSS VSS VCC VCC _2442_ sky130_fd_sc_hs__mux2_1
X_4045_ _1665_ _1686_ _1688_ VSS VSS VCC VCC _0077_ sky130_fd_sc_hs__a21o_1
X_4947_ _2304_ _2306_ VSS VSS VCC VCC _2307_ sky130_fd_sc_hs__xnor2_1
X_4878_ u_muldiv.o_div\[29\] _2264_ u_muldiv.o_div\[30\] VSS VSS VCC VCC _2272_
+ sky130_fd_sc_hs__o21ai_1
X_3829_ _0628_ _1542_ _1545_ _1548_ VSS VSS VCC VCC _1549_ sky130_fd_sc_hs__or4_1
Xclkbuf_leaf_40_i_clk clknet_2_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_40_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_4801_ u_muldiv.quotient_msk\[14\] u_muldiv.o_div\[14\] _1841_ VSS VSS VCC
+ VCC _2211_ sky130_fd_sc_hs__o21a_1
X_5781_ clknet_leaf_28_i_clk _0423_ VSS VSS VCC VCC u_muldiv.o_div\[0\] sky130_fd_sc_hs__dfxtp_1
X_2993_ _0746_ _0805_ _0447_ VSS VSS VCC VCC _0806_ sky130_fd_sc_hs__a21o_1
X_4732_ u_muldiv.o_div\[1\] _2029_ _2154_ VSS VSS VCC VCC _2155_ sky130_fd_sc_hs__mux2_1
X_4663_ _2084_ _2085_ VSS VSS VCC VCC _2086_ sky130_fd_sc_hs__nand2_1
X_3614_ _0670_ _0794_ _0867_ VSS VSS VCC VCC _1348_ sky130_fd_sc_hs__a21o_1
X_4594_ _1204_ _2019_ _2020_ VSS VSS VCC VCC _0294_ sky130_fd_sc_hs__nor3_1
X_3545_ _1250_ u_bits.i_op1\[10\] _1251_ _0777_ _0778_ _0783_ VSS VSS VCC VCC
+ _1281_ sky130_fd_sc_hs__mux4_1
X_3476_ o_wdata[4] u_wr_mux.i_reg_data2\[20\] _1224_ VSS VSS VCC VCC _1229_
+ sky130_fd_sc_hs__mux2_1
X_5215_ u_muldiv.dividend\[25\] u_muldiv.dividend\[24\] _2525_ VSS VSS VCC VCC
+ _2552_ sky130_fd_sc_hs__or3_2
X_5146_ _2084_ _2479_ VSS VSS VCC VCC _2489_ sky130_fd_sc_hs__nand2_1
X_5077_ _2044_ _2415_ _2425_ VSS VSS VCC VCC _2426_ sky130_fd_sc_hs__a21oi_1
X_4028_ _1665_ _1674_ _1676_ VSS VSS VCC VCC _0072_ sky130_fd_sc_hs__a21o_1
X_3330_ _1108_ _1122_ _0446_ VSS VSS VCC VCC _1123_ sky130_fd_sc_hs__a21o_1
X_5000_ _2355_ VSS VSS VCC VCC _0365_ sky130_fd_sc_hs__clkbuf_1
X_3261_ _0775_ _1057_ _0784_ _0945_ _0879_ _0789_ VSS VSS VCC VCC _1058_ sky130_fd_sc_hs__mux4_2
X_3192_ _0993_ VSS VSS VCC VCC o_add[27] sky130_fd_sc_hs__inv_2
X_5764_ clknet_leaf_18_i_clk _0407_ VSS VSS VCC VCC u_muldiv.divisor\[16\]
+ sky130_fd_sc_hs__dfxtp_1
X_2976_ _0758_ VSS VSS VCC VCC _0789_ sky130_fd_sc_hs__buf_4
X_5695_ clknet_leaf_29_i_clk _0338_ VSS VSS VCC VCC u_muldiv.quotient_msk\[9\]
+ sky130_fd_sc_hs__dfxtp_1
X_4715_ _2136_ u_muldiv.dividend\[30\] _2137_ VSS VSS VCC VCC _2138_ sky130_fd_sc_hs__a21o_1
X_4646_ _2058_ _2067_ _2068_ VSS VSS VCC VCC _2069_ sky130_fd_sc_hs__a21boi_1
X_4577_ o_add[25] _2004_ VSS VSS VCC VCC _2013_ sky130_fd_sc_hs__and2_1
X_3528_ _0642_ _0683_ VSS VSS VCC VCC _1265_ sky130_fd_sc_hs__or2_2
X_3459_ u_wr_mux.i_reg_data2\[12\] o_wdata[4] _0718_ VSS VSS VCC VCC _1220_
+ sky130_fd_sc_hs__mux2_1
X_5129_ _1841_ _2466_ _2473_ VSS VSS VCC VCC _2474_ sky130_fd_sc_hs__a21o_1
X_2830_ u_bits.i_op1\[18\] VSS VSS VCC VCC _0645_ sky130_fd_sc_hs__buf_4
X_2761_ _0569_ _0570_ _0562_ _0574_ _0575_ VSS VSS VCC VCC _0576_ sky130_fd_sc_hs__o221a_2
X_4500_ _1981_ VSS VSS VCC VCC _0239_ sky130_fd_sc_hs__clkbuf_1
X_2692_ _0505_ _0506_ VSS VSS VCC VCC _0507_ sky130_fd_sc_hs__nand2_1
X_5480_ clknet_leaf_1_i_clk _0128_ VSS VSS VCC VCC u_bits.i_sra sky130_fd_sc_hs__dfxtp_2
X_4431_ u_muldiv.divisor\[52\] _1836_ _1887_ u_muldiv.divisor\[53\] _1933_ VSS VSS
+ VCC VCC _0218_ sky130_fd_sc_hs__a221o_1
X_4362_ _1877_ VSS VSS VCC VCC _1878_ sky130_fd_sc_hs__buf_4
X_4293_ _1821_ VSS VSS VCC VCC _0192_ sky130_fd_sc_hs__clkbuf_1
X_3313_ _0728_ VSS VSS VCC VCC _1106_ sky130_fd_sc_hs__buf_2
X_3244_ _0461_ u_bits.i_op2\[29\] _0465_ u_bits.i_op1\[29\] VSS VSS VCC VCC
+ _1042_ sky130_fd_sc_hs__a22o_1
X_3175_ _0689_ u_bits.i_op2\[26\] VSS VSS VCC VCC _0978_ sky130_fd_sc_hs__nand2_1
X_5747_ clknet_leaf_21_i_clk _0390_ VSS VSS VCC VCC u_muldiv.dividend\[31\]
+ sky130_fd_sc_hs__dfxtp_2
X_2959_ u_bits.i_op1\[21\] _0630_ _0656_ VSS VSS VCC VCC _0772_ sky130_fd_sc_hs__mux2_1
X_5678_ clknet_leaf_31_i_clk _0321_ VSS VSS VCC VCC u_muldiv.o_div\[24\] sky130_fd_sc_hs__dfxtp_1
X_4629_ u_muldiv.divisor\[8\] u_muldiv.dividend\[8\] VSS VSS VCC VCC _2052_
+ sky130_fd_sc_hs__or2b_1
X_4980_ _2070_ _2057_ _2069_ VSS VSS VCC VCC _2337_ sky130_fd_sc_hs__o21a_1
X_3931_ _1617_ VSS VSS VCC VCC _0034_ sky130_fd_sc_hs__clkbuf_1
X_3862_ _1214_ VSS VSS VCC VCC _1579_ sky130_fd_sc_hs__clkbuf_2
X_5601_ clknet_leaf_32_i_clk _0248_ VSS VSS VCC VCC u_muldiv.mul\[18\] sky130_fd_sc_hs__dfxtp_1
X_2813_ _0627_ VSS VSS VCC VCC _0628_ sky130_fd_sc_hs__buf_2
X_5532_ clknet_leaf_14_i_clk _0180_ VSS VSS VCC VCC csr_data\[16\] sky130_fd_sc_hs__dfxtp_1
X_3793_ u_bits.i_op2\[15\] _0654_ _1267_ VSS VSS VCC VCC _1515_ sky130_fd_sc_hs__a21oi_1
X_2744_ _0455_ _0558_ VSS VSS VCC VCC _0559_ sky130_fd_sc_hs__xnor2_4
X_5463_ clknet_leaf_10_i_clk _0111_ VSS VSS VCC VCC o_pc_target[5] sky130_fd_sc_hs__dfxtp_2
X_2675_ _0457_ _0489_ VSS VSS VCC VCC _0490_ sky130_fd_sc_hs__xnor2_1
X_5394_ clknet_leaf_53_i_clk _0042_ VSS VSS VCC VCC u_bits.i_op1\[26\] sky130_fd_sc_hs__dfxtp_2
X_4414_ _1850_ _1919_ VSS VSS VCC VCC _1920_ sky130_fd_sc_hs__nand2_1
X_4345_ _1376_ _1863_ VSS VSS VCC VCC _1864_ sky130_fd_sc_hs__nand2_1
X_4276_ csr_data\[20\] i_csr_data[20] _1811_ VSS VSS VCC VCC _1813_ sky130_fd_sc_hs__mux2_1
X_3227_ u_muldiv.mul\[28\] _0740_ _0720_ u_muldiv.mul\[60\] _1025_ VSS VSS VCC
+ VCC _1026_ sky130_fd_sc_hs__a221o_1
X_3158_ _0960_ _0961_ VSS VSS VCC VCC _0962_ sky130_fd_sc_hs__nand2_1
X_3089_ _0461_ u_bits.i_op2\[24\] _0465_ u_bits.i_op1\[24\] VSS VSS VCC VCC
+ _0897_ sky130_fd_sc_hs__a22o_1
X_4130_ o_pc_target[8] i_pc_target[8] _1734_ VSS VSS VCC VCC _1737_ sky130_fd_sc_hs__mux2_1
X_4061_ _1689_ _1698_ _1699_ VSS VSS VCC VCC _0082_ sky130_fd_sc_hs__a21o_1
X_3012_ _0779_ _0700_ _0762_ VSS VSS VCC VCC _0823_ sky130_fd_sc_hs__o21a_1
X_4963_ _0794_ _2321_ VSS VSS VCC VCC _2322_ sky130_fd_sc_hs__xor2_1
X_3914_ _1608_ VSS VSS VCC VCC _0026_ sky130_fd_sc_hs__clkbuf_1
X_4894_ u_muldiv.quotient_msk\[6\] _1210_ _2279_ u_muldiv.quotient_msk\[7\] VSS
+ VSS VCC VCC _0335_ sky130_fd_sc_hs__a22o_1
X_3845_ _0749_ o_add[18] _1562_ _1563_ _0453_ VSS VSS VCC VCC _1564_ sky130_fd_sc_hs__a221o_1
X_3776_ _0818_ _0822_ _1309_ _1314_ _0758_ _0673_ VSS VSS VCC VCC _1499_ sky130_fd_sc_hs__mux4_1
X_5515_ clknet_leaf_10_i_clk _0163_ VSS VSS VCC VCC o_to_trap sky130_fd_sc_hs__dfxtp_2
X_2727_ _0539_ _0540_ _0541_ VSS VSS VCC VCC _0542_ sky130_fd_sc_hs__mux2_2
X_5446_ clknet_leaf_9_i_clk _0094_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[6\]
+ sky130_fd_sc_hs__dfxtp_1
X_2658_ u_bits.i_op1\[19\] u_muldiv.add_prev\[19\] _0451_ VSS VSS VCC VCC
+ _0473_ sky130_fd_sc_hs__mux2_1
X_5377_ clknet_leaf_47_i_clk _0025_ VSS VSS VCC VCC u_bits.i_op1\[9\] sky130_fd_sc_hs__dfxtp_2
X_4328_ _1845_ VSS VSS VCC VCC _1850_ sky130_fd_sc_hs__buf_2
X_4259_ csr_data\[12\] i_csr_data[12] _1800_ VSS VSS VCC VCC _1804_ sky130_fd_sc_hs__mux2_1
X_3630_ _0687_ _1310_ _1267_ VSS VSS VCC VCC _1363_ sky130_fd_sc_hs__a21oi_1
X_3561_ _1249_ _1291_ _1296_ VSS VSS VCC VCC _1297_ sky130_fd_sc_hs__a21bo_1
X_5300_ u_muldiv.divisor\[14\] _2614_ _2615_ u_muldiv.divisor\[15\] VSS VSS VCC
+ VCC _0405_ sky130_fd_sc_hs__a22o_1
X_3492_ _1192_ u_wr_mux.i_reg_data2\[27\] _1237_ VSS VSS VCC VCC o_wdata[27]
+ sky130_fd_sc_hs__a21o_2
X_5231_ _2117_ _2557_ _2114_ VSS VSS VCC VCC _2566_ sky130_fd_sc_hs__a21oi_1
X_5162_ _2498_ _2503_ _1877_ VSS VSS VCC VCC _2504_ sky130_fd_sc_hs__mux2_1
X_5093_ _2436_ _2438_ _2440_ _2375_ VSS VSS VCC VCC _2441_ sky130_fd_sc_hs__a22o_1
X_4113_ i_res_src[1] _1638_ _1635_ _0730_ VSS VSS VCC VCC _0105_ sky130_fd_sc_hs__a22o_1
X_4044_ u_bits.i_op2\[20\] _1687_ _1675_ i_op2[20] VSS VSS VCC VCC _1688_
+ sky130_fd_sc_hs__a22o_1
X_4946_ _2061_ _2305_ VSS VSS VCC VCC _2306_ sky130_fd_sc_hs__nand2_1
X_4877_ u_muldiv.o_div\[29\] u_muldiv.o_div\[30\] _2264_ _1207_ VSS VSS VCC
+ VCC _2271_ sky130_fd_sc_hs__o31a_1
X_3828_ _0672_ _1546_ _1547_ _0800_ VSS VSS VCC VCC _1548_ sky130_fd_sc_hs__o211a_1
X_3759_ _1333_ csr_data\[12\] _1388_ VSS VSS VCC VCC _1484_ sky130_fd_sc_hs__o21ai_1
X_5429_ clknet_leaf_1_i_clk _0077_ VSS VSS VCC VCC u_bits.i_op2\[20\] sky130_fd_sc_hs__dfxtp_4
X_4800_ u_muldiv.o_div\[13\] u_muldiv.o_div\[14\] _2201_ VSS VSS VCC VCC _2210_
+ sky130_fd_sc_hs__or3_2
X_2992_ _0750_ o_add[21] _0802_ _0803_ _0804_ VSS VSS VCC VCC _0805_ sky130_fd_sc_hs__a221o_1
X_5780_ clknet_leaf_5_i_clk _0003_ VSS VSS VCC VCC u_muldiv.add_prev\[31\]
+ sky130_fd_sc_hs__dfxtp_1
X_4731_ _2153_ VSS VSS VCC VCC _2154_ sky130_fd_sc_hs__buf_4
X_4662_ u_muldiv.dividend\[18\] u_muldiv.divisor\[18\] VSS VSS VCC VCC _2085_
+ sky130_fd_sc_hs__or2b_1
X_3613_ _0669_ _0788_ _0881_ VSS VSS VCC VCC _1347_ sky130_fd_sc_hs__or3b_1
X_4593_ op_cnt\[0\] op_cnt\[1\] op_cnt\[2\] VSS VSS VCC VCC _2020_ sky130_fd_sc_hs__and3_1
X_3544_ _0447_ _1279_ _1280_ _1124_ VSS VSS VCC VCC o_result[0] sky130_fd_sc_hs__o211a_2
X_3475_ _1228_ VSS VSS VCC VCC o_wdata[19] sky130_fd_sc_hs__buf_2
X_5214_ u_muldiv.dividend\[24\] _2525_ u_muldiv.dividend\[25\] VSS VSS VCC VCC
+ _2551_ sky130_fd_sc_hs__o21ai_1
X_5145_ u_muldiv.dividend\[18\] _2468_ u_muldiv.dividend\[19\] VSS VSS VCC VCC
+ _2488_ sky130_fd_sc_hs__o21ai_1
X_5076_ _2043_ _2080_ VSS VSS VCC VCC _2425_ sky130_fd_sc_hs__and2b_1
X_4027_ u_bits.i_op2\[15\] _1663_ _1675_ i_op2[15] VSS VSS VCC VCC _1676_
+ sky130_fd_sc_hs__a22o_1
X_4929_ _2062_ _2063_ VSS VSS VCC VCC _2290_ sky130_fd_sc_hs__nor2_1
X_3260_ _1056_ _1001_ _0774_ VSS VSS VCC VCC _1057_ sky130_fd_sc_hs__mux2_1
X_3191_ _0991_ _0992_ VSS VSS VCC VCC _0993_ sky130_fd_sc_hs__xnor2_2
X_5763_ clknet_leaf_19_i_clk _0406_ VSS VSS VCC VCC u_muldiv.divisor\[15\]
+ sky130_fd_sc_hs__dfxtp_1
X_4714_ _1834_ u_muldiv.dividend\[31\] VSS VSS VCC VCC _2137_ sky130_fd_sc_hs__and2_1
X_2975_ _0524_ VSS VSS VCC VCC _0788_ sky130_fd_sc_hs__clkbuf_4
X_5694_ clknet_leaf_27_i_clk _0337_ VSS VSS VCC VCC u_muldiv.quotient_msk\[8\]
+ sky130_fd_sc_hs__dfxtp_1
X_4645_ u_muldiv.divisor\[4\] u_muldiv.dividend\[4\] VSS VSS VCC VCC _2068_
+ sky130_fd_sc_hs__or2b_1
X_4576_ _0903_ _2007_ VSS VSS VCC VCC _0284_ sky130_fd_sc_hs__nor2_1
X_3527_ _1249_ _1263_ VSS VSS VCC VCC _1264_ sky130_fd_sc_hs__nand2_1
X_3458_ _1219_ VSS VSS VCC VCC o_wdata[11] sky130_fd_sc_hs__buf_2
X_3389_ _0480_ _1166_ VSS VSS VCC VCC o_add[19] sky130_fd_sc_hs__xnor2_4
X_5128_ _1207_ _2467_ _2468_ _2472_ VSS VSS VCC VCC _2473_ sky130_fd_sc_hs__a31o_1
X_5059_ _1251_ _2409_ VSS VSS VCC VCC _2410_ sky130_fd_sc_hs__xnor2_1
X_2760_ _0554_ _0555_ VSS VSS VCC VCC _0575_ sky130_fd_sc_hs__nand2_1
X_2691_ u_bits.i_op1\[14\] u_muldiv.add_prev\[14\] _0449_ VSS VSS VCC VCC
+ _0506_ sky130_fd_sc_hs__mux2_2
X_4430_ _1832_ _1932_ VSS VSS VCC VCC _1933_ sky130_fd_sc_hs__nor2_1
X_4361_ _1827_ VSS VSS VCC VCC _1877_ sky130_fd_sc_hs__clkbuf_4
X_4292_ csr_data\[28\] i_csr_data[28] _1811_ VSS VSS VCC VCC _1821_ sky130_fd_sc_hs__mux2_1
X_3312_ _1104_ _1105_ VSS VSS VCC VCC o_add[31] sky130_fd_sc_hs__nor2_4
X_3243_ _0739_ csr_data\[28\] _1041_ _0732_ VSS VSS VCC VCC o_result[28] sky130_fd_sc_hs__o211a_2
X_3174_ _0833_ _0976_ _0835_ _0832_ _0879_ _0789_ VSS VSS VCC VCC _0977_ sky130_fd_sc_hs__mux4_1
X_5746_ clknet_leaf_22_i_clk _0389_ VSS VSS VCC VCC u_muldiv.dividend\[30\]
+ sky130_fd_sc_hs__dfxtp_4
X_2958_ _0768_ u_bits.i_op2\[21\] _0637_ _0770_ VSS VSS VCC VCC _0771_ sky130_fd_sc_hs__o22a_1
X_5677_ clknet_leaf_31_i_clk _0320_ VSS VSS VCC VCC u_muldiv.o_div\[23\] sky130_fd_sc_hs__dfxtp_1
X_4628_ u_muldiv.dividend\[9\] u_muldiv.divisor\[9\] VSS VSS VCC VCC _2051_
+ sky130_fd_sc_hs__and2b_1
X_2889_ u_bits.i_op2\[2\] _0703_ VSS VSS VCC VCC _0704_ sky130_fd_sc_hs__nand2_1
X_4559_ _1157_ _2007_ VSS VSS VCC VCC _0272_ sky130_fd_sc_hs__nor2_1
X_3930_ _0645_ i_op1[18] _1610_ VSS VSS VCC VCC _1617_ sky130_fd_sc_hs__mux2_1
X_3861_ _1106_ csr_data\[19\] _1578_ _1124_ VSS VSS VCC VCC o_result[19] sky130_fd_sc_hs__o211a_2
X_5600_ clknet_leaf_32_i_clk _0247_ VSS VSS VCC VCC u_muldiv.mul\[17\] sky130_fd_sc_hs__dfxtp_1
X_3792_ _0688_ _1512_ _1513_ _1249_ VSS VSS VCC VCC _1514_ sky130_fd_sc_hs__o211a_1
X_2812_ _0625_ _0626_ VSS VSS VCC VCC _0627_ sky130_fd_sc_hs__nor2_1
X_5531_ clknet_leaf_14_i_clk _0179_ VSS VSS VCC VCC csr_data\[15\] sky130_fd_sc_hs__dfxtp_1
X_2743_ _0448_ u_bits.i_op1\[6\] _0497_ _0557_ VSS VSS VCC VCC _0558_ sky130_fd_sc_hs__a31o_1
X_5462_ clknet_leaf_10_i_clk _0110_ VSS VSS VCC VCC o_pc_target[4] sky130_fd_sc_hs__dfxtp_2
X_2674_ _0460_ u_bits.i_op2\[16\] u_bits.i_op1\[16\] _0464_ VSS VSS VCC VCC
+ _0489_ sky130_fd_sc_hs__a22o_1
X_5393_ clknet_leaf_53_i_clk _0041_ VSS VSS VCC VCC u_bits.i_op1\[25\] sky130_fd_sc_hs__dfxtp_2
X_4413_ u_bits.i_op2\[16\] u_bits.i_op2\[17\] _1910_ VSS VSS VCC VCC _1919_
+ sky130_fd_sc_hs__or3_1
X_4344_ _0688_ _1859_ _1846_ VSS VSS VCC VCC _1863_ sky130_fd_sc_hs__o21ai_1
X_4275_ _1812_ VSS VSS VCC VCC _0183_ sky130_fd_sc_hs__clkbuf_1
X_3226_ u_muldiv.dividend\[28\] _0721_ _0723_ u_muldiv.o_div\[28\] _0744_ VSS VSS
+ VCC VCC _1025_ sky130_fd_sc_hs__a221o_1
X_3157_ u_bits.i_op1\[26\] u_muldiv.add_prev\[26\] _0451_ VSS VSS VCC VCC
+ _0961_ sky130_fd_sc_hs__mux2_1
X_3088_ _0496_ _0614_ _0736_ _0893_ _0469_ VSS VSS VCC VCC _0896_ sky130_fd_sc_hs__a2111o_1
X_5729_ clknet_leaf_19_i_clk _0372_ VSS VSS VCC VCC u_muldiv.dividend\[13\]
+ sky130_fd_sc_hs__dfxtp_2
X_4060_ u_bits.i_op2\[25\] _1687_ _1596_ i_op2[25] VSS VSS VCC VCC _1699_
+ sky130_fd_sc_hs__a22o_1
X_3011_ _0821_ VSS VSS VCC VCC _0822_ sky130_fd_sc_hs__inv_2
X_4962_ _1255_ _2308_ _2292_ VSS VSS VCC VCC _2321_ sky130_fd_sc_hs__o21a_1
X_4893_ u_muldiv.quotient_msk\[5\] _1210_ _2279_ u_muldiv.quotient_msk\[6\] VSS
+ VSS VCC VCC _0334_ sky130_fd_sc_hs__a22o_1
X_3913_ _1305_ i_op1[10] _1599_ VSS VSS VCC VCC _1608_ sky130_fd_sc_hs__mux2_1
X_3844_ _0908_ _1556_ _0955_ VSS VSS VCC VCC _1563_ sky130_fd_sc_hs__a21oi_1
X_3775_ _1497_ _1498_ _0730_ u_pc_sel.i_pc_next\[13\] VSS VSS VCC VCC o_result[13]
+ sky130_fd_sc_hs__a2bb2o_2
X_5514_ clknet_leaf_12_i_clk _0162_ VSS VSS VCC VCC csr_read sky130_fd_sc_hs__dfxtp_1
X_2726_ _0459_ u_bits.i_op2\[0\] u_bits.i_op1\[0\] _0463_ VSS VSS VCC VCC
+ _0541_ sky130_fd_sc_hs__a22o_2
X_2657_ _0457_ _0471_ VSS VSS VCC VCC _0472_ sky130_fd_sc_hs__xnor2_1
X_5445_ clknet_leaf_2_i_clk _0093_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[5\]
+ sky130_fd_sc_hs__dfxtp_1
X_5376_ clknet_leaf_47_i_clk _0024_ VSS VSS VCC VCC u_bits.i_op1\[8\] sky130_fd_sc_hs__dfxtp_2
X_4327_ u_muldiv.divisor\[32\] _1838_ _1843_ u_muldiv.divisor\[33\] _1849_ VSS VSS
+ VCC VCC _0198_ sky130_fd_sc_hs__a221o_1
X_4258_ _1803_ VSS VSS VCC VCC _0175_ sky130_fd_sc_hs__clkbuf_1
X_3209_ _0628_ _1000_ _1009_ _0747_ VSS VSS VCC VCC _1010_ sky130_fd_sc_hs__o31a_1
X_4189_ u_wr_mux.i_reg_data2\[12\] i_reg_data2[12] _1767_ VSS VSS VCC VCC
+ _1768_ sky130_fd_sc_hs__mux2_1
X_3560_ _1265_ _1292_ _1295_ _0634_ VSS VSS VCC VCC _1296_ sky130_fd_sc_hs__o211a_1
X_5230_ u_muldiv.dividend\[26\] _2552_ u_muldiv.dividend\[27\] VSS VSS VCC VCC
+ _2565_ sky130_fd_sc_hs__o21ai_1
X_3491_ o_wdata[3] _1233_ _0799_ u_wr_mux.i_reg_data2\[11\] VSS VSS VCC VCC
+ _1237_ sky130_fd_sc_hs__a22o_1
X_5161_ _2500_ _2502_ _2288_ VSS VSS VCC VCC _2503_ sky130_fd_sc_hs__mux2_1
X_5092_ _0655_ _2439_ VSS VSS VCC VCC _2440_ sky130_fd_sc_hs__xnor2_1
X_4112_ i_res_src[0] _1638_ _1636_ o_res_src[0] VSS VSS VCC VCC _0104_ sky130_fd_sc_hs__a22o_1
X_4043_ _1634_ VSS VSS VCC VCC _1687_ sky130_fd_sc_hs__buf_2
X_4945_ _2060_ u_muldiv.dividend\[2\] VSS VSS VCC VCC _2305_ sky130_fd_sc_hs__nand2_1
X_4876_ _2167_ _2268_ _2270_ VSS VSS VCC VCC _0326_ sky130_fd_sc_hs__a21oi_1
X_3827_ _0687_ _1292_ VSS VSS VCC VCC _1547_ sky130_fd_sc_hs__nand2_1
X_3758_ _1331_ _1479_ _1481_ _1482_ _1357_ VSS VSS VCC VCC _1483_ sky130_fd_sc_hs__o221a_1
X_2709_ u_bits.i_op2\[3\] VSS VSS VCC VCC _0524_ sky130_fd_sc_hs__buf_4
X_3689_ _1254_ _1262_ _0910_ _0824_ _0670_ _0643_ VSS VSS VCC VCC _1418_ sky130_fd_sc_hs__mux4_1
X_5428_ clknet_leaf_52_i_clk _0076_ VSS VSS VCC VCC u_bits.i_op2\[19\] sky130_fd_sc_hs__dfxtp_4
X_5359_ clknet_leaf_40_i_clk _0007_ VSS VSS VCC VCC u_muldiv.mul\[55\] sky130_fd_sc_hs__dfxtp_1
X_2991_ _0452_ VSS VSS VCC VCC _0804_ sky130_fd_sc_hs__clkbuf_4
X_4730_ u_muldiv.outsign _1206_ _2152_ VSS VSS VCC VCC _2153_ sky130_fd_sc_hs__a21o_2
X_4661_ u_muldiv.divisor\[18\] u_muldiv.dividend\[18\] VSS VSS VCC VCC _2084_
+ sky130_fd_sc_hs__or2b_1
X_3612_ _1342_ _1345_ _0644_ VSS VSS VCC VCC _1346_ sky130_fd_sc_hs__mux2_1
X_4592_ op_cnt\[0\] op_cnt\[1\] op_cnt\[2\] VSS VSS VCC VCC _2019_ sky130_fd_sc_hs__a21oi_1
X_3543_ _0728_ csr_data\[0\] VSS VSS VCC VCC _1280_ sky130_fd_sc_hs__or2_1
X_3474_ o_wdata[3] u_wr_mux.i_reg_data2\[19\] _1224_ VSS VSS VCC VCC _1228_
+ sky130_fd_sc_hs__mux2_1
X_5213_ _2362_ _2548_ _0943_ VSS VSS VCC VCC _2550_ sky130_fd_sc_hs__a21oi_1
X_5144_ u_muldiv.dividend\[19\] u_muldiv.dividend\[18\] _2468_ VSS VSS VCC VCC
+ _2487_ sky130_fd_sc_hs__or3_1
X_5075_ u_muldiv.dividend\[12\] _2403_ u_muldiv.dividend\[13\] VSS VSS VCC VCC
+ _2424_ sky130_fd_sc_hs__o21ai_1
X_4026_ _1595_ VSS VSS VCC VCC _1675_ sky130_fd_sc_hs__buf_2
X_4928_ _2062_ _2063_ VSS VSS VCC VCC _2289_ sky130_fd_sc_hs__and2_1
X_4859_ u_muldiv.o_div\[25\] _2250_ u_muldiv.o_div\[26\] VSS VSS VCC VCC _2257_
+ sky130_fd_sc_hs__o21ai_1
X_3190_ _0964_ _0967_ _0962_ VSS VSS VCC VCC _0992_ sky130_fd_sc_hs__a21bo_1
X_5762_ clknet_leaf_19_i_clk _0405_ VSS VSS VCC VCC u_muldiv.divisor\[14\]
+ sky130_fd_sc_hs__dfxtp_1
X_2974_ u_bits.i_op1\[9\] _0785_ u_bits.i_op1\[7\] _0786_ _0658_ _0659_ VSS VSS
+ VCC VCC _0787_ sky130_fd_sc_hs__mux4_2
X_4713_ u_muldiv.divisor\[30\] VSS VSS VCC VCC _2136_ sky130_fd_sc_hs__inv_2
X_5693_ clknet_leaf_27_i_clk _0336_ VSS VSS VCC VCC u_muldiv.quotient_msk\[7\]
+ sky130_fd_sc_hs__dfxtp_1
X_4644_ _2059_ _2061_ _2065_ _2066_ VSS VSS VCC VCC _2067_ sky130_fd_sc_hs__a31o_1
X_4575_ _0855_ _2007_ VSS VSS VCC VCC _0283_ sky130_fd_sc_hs__nor2_1
X_3526_ _1254_ _1260_ _0910_ _1262_ _0674_ _0644_ VSS VSS VCC VCC _1263_ sky130_fd_sc_hs__mux4_1
X_3457_ u_wr_mux.i_reg_data2\[11\] o_wdata[3] _0718_ VSS VSS VCC VCC _1219_
+ sky130_fd_sc_hs__mux2_1
X_3388_ _0482_ _1165_ _0478_ VSS VSS VCC VCC _1166_ sky130_fd_sc_hs__o21a_1
X_5127_ _1880_ _2470_ _2471_ VSS VSS VCC VCC _2472_ sky130_fd_sc_hs__and3_1
X_5058_ _1305_ _2394_ _2293_ VSS VSS VCC VCC _2409_ sky130_fd_sc_hs__o21a_1
X_4009_ _1634_ VSS VSS VCC VCC _1663_ sky130_fd_sc_hs__buf_2
X_2690_ _0456_ _0504_ VSS VSS VCC VCC _0505_ sky130_fd_sc_hs__xnor2_4
X_4360_ u_muldiv.divisor\[38\] _1867_ _1843_ u_muldiv.divisor\[39\] _1876_ VSS VSS
+ VCC VCC _0204_ sky130_fd_sc_hs__a221o_1
X_3311_ _1070_ _1094_ _1103_ VSS VSS VCC VCC _1105_ sky130_fd_sc_hs__and3_1
X_4291_ _1820_ VSS VSS VCC VCC _0191_ sky130_fd_sc_hs__clkbuf_1
X_3242_ _1026_ _1040_ _0447_ VSS VSS VCC VCC _1041_ sky130_fd_sc_hs__a21o_1
X_3173_ _0689_ _0943_ _0904_ _0692_ _0651_ _0774_ VSS VSS VCC VCC _0976_ sky130_fd_sc_hs__mux4_1
X_5745_ clknet_leaf_21_i_clk _0388_ VSS VSS VCC VCC u_muldiv.dividend\[29\]
+ sky130_fd_sc_hs__dfxtp_2
X_2957_ _0618_ _0639_ _0769_ VSS VSS VCC VCC _0770_ sky130_fd_sc_hs__and3_1
X_5676_ clknet_leaf_30_i_clk _0319_ VSS VSS VCC VCC u_muldiv.o_div\[22\] sky130_fd_sc_hs__dfxtp_1
X_2888_ _0702_ u_bits.i_sra VSS VSS VCC VCC _0703_ sky130_fd_sc_hs__nand2_4
X_4627_ _2048_ _2049_ VSS VSS VCC VCC _2050_ sky130_fd_sc_hs__nand2_1
X_4558_ _1214_ VSS VSS VCC VCC _2007_ sky130_fd_sc_hs__clkbuf_4
X_4489_ _1975_ VSS VSS VCC VCC _0234_ sky130_fd_sc_hs__clkbuf_1
X_3509_ _0620_ _1195_ VSS VSS VCC VCC _1246_ sky130_fd_sc_hs__nand2_1
Xclkbuf_2_3__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_3__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_3860_ _1567_ _1577_ _0446_ VSS VSS VCC VCC _1578_ sky130_fd_sc_hs__a21o_1
X_3791_ _0860_ _0911_ _0687_ VSS VSS VCC VCC _1513_ sky130_fd_sc_hs__a21bo_1
X_2811_ o_funct3[1] o_funct3[0] VSS VSS VCC VCC _0626_ sky130_fd_sc_hs__nand2_2
X_5530_ clknet_leaf_14_i_clk _0178_ VSS VSS VCC VCC csr_data\[14\] sky130_fd_sc_hs__dfxtp_1
X_2742_ u_mux.i_group_mux u_bits.i_op2\[6\] VSS VSS VCC VCC _0557_ sky130_fd_sc_hs__and2b_1
Xclkbuf_leaf_53_i_clk clknet_2_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_53_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_5461_ clknet_leaf_13_i_clk _0109_ VSS VSS VCC VCC o_pc_target[3] sky130_fd_sc_hs__dfxtp_2
X_2673_ _0486_ _0487_ VSS VSS VCC VCC _0488_ sky130_fd_sc_hs__nand2_1
X_4412_ u_muldiv.divisor\[48\] _1867_ _1887_ u_muldiv.divisor\[49\] _1918_ VSS VSS
+ VCC VCC _0214_ sky130_fd_sc_hs__a221o_1
X_5392_ clknet_leaf_53_i_clk _0040_ VSS VSS VCC VCC u_bits.i_op1\[24\] sky130_fd_sc_hs__dfxtp_2
X_4343_ u_muldiv.divisor\[35\] _1838_ _1843_ u_muldiv.divisor\[36\] _1862_ VSS VSS
+ VCC VCC _0201_ sky130_fd_sc_hs__a221o_1
X_4274_ csr_data\[19\] i_csr_data[19] _1811_ VSS VSS VCC VCC _1812_ sky130_fd_sc_hs__mux2_1
X_3225_ _1024_ VSS VSS VCC VCC o_add[28] sky130_fd_sc_hs__inv_2
X_3156_ _0458_ _0959_ VSS VSS VCC VCC _0960_ sky130_fd_sc_hs__xnor2_1
X_3087_ _0810_ _0852_ _0893_ _0814_ _0894_ VSS VSS VCC VCC _0895_ sky130_fd_sc_hs__o221a_1
X_5728_ clknet_leaf_20_i_clk _0371_ VSS VSS VCC VCC u_muldiv.dividend\[12\]
+ sky130_fd_sc_hs__dfxtp_2
X_3989_ _0688_ _1637_ _1638_ i_op2[4] VSS VSS VCC VCC _1649_ sky130_fd_sc_hs__a22o_1
X_5659_ clknet_leaf_27_i_clk _0302_ VSS VSS VCC VCC u_muldiv.o_div\[5\] sky130_fd_sc_hs__dfxtp_1
X_3010_ _0648_ _0698_ _0820_ VSS VSS VCC VCC _0821_ sky130_fd_sc_hs__a21oi_1
X_4961_ _2061_ _2065_ _2318_ _1839_ VSS VSS VCC VCC _2320_ sky130_fd_sc_hs__a31o_1
X_4892_ u_muldiv.quotient_msk\[4\] _1210_ _2279_ u_muldiv.quotient_msk\[5\] VSS
+ VSS VCC VCC _0333_ sky130_fd_sc_hs__a22o_1
X_3912_ _1607_ VSS VSS VCC VCC _0025_ sky130_fd_sc_hs__clkbuf_1
X_3843_ _0858_ _1555_ _1558_ _1561_ VSS VSS VCC VCC _1562_ sky130_fd_sc_hs__or4_1
X_3774_ _1333_ csr_data\[13\] _1388_ VSS VSS VCC VCC _1498_ sky130_fd_sc_hs__o21ai_1
X_5513_ clknet_leaf_47_i_clk _0161_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[31\]
+ sky130_fd_sc_hs__dfxtp_2
X_2725_ u_bits.i_op1\[0\] u_muldiv.add_prev\[0\] _0449_ VSS VSS VCC VCC _0540_
+ sky130_fd_sc_hs__mux2_2
X_2656_ _0460_ u_bits.i_op2\[19\] u_bits.i_op1\[19\] _0464_ VSS VSS VCC VCC
+ _0471_ sky130_fd_sc_hs__a22o_1
X_5444_ clknet_leaf_2_i_clk _0092_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[4\]
+ sky130_fd_sc_hs__dfxtp_1
X_5375_ clknet_leaf_47_i_clk _0023_ VSS VSS VCC VCC u_bits.i_op1\[7\] sky130_fd_sc_hs__dfxtp_2
X_4326_ _1832_ _1848_ VSS VSS VCC VCC _1849_ sky130_fd_sc_hs__nor2_1
X_4257_ csr_data\[11\] i_csr_data[11] _1800_ VSS VSS VCC VCC _1803_ sky130_fd_sc_hs__mux2_1
X_4188_ _1711_ VSS VSS VCC VCC _1767_ sky130_fd_sc_hs__clkbuf_4
X_3208_ _0925_ _1003_ _1006_ _0914_ _1008_ VSS VSS VCC VCC _1009_ sky130_fd_sc_hs__a221o_1
X_3139_ _0943_ _0904_ _0658_ VSS VSS VCC VCC _0944_ sky130_fd_sc_hs__mux2_1
X_3490_ _1192_ u_wr_mux.i_reg_data2\[26\] _1236_ VSS VSS VCC VCC o_wdata[26]
+ sky130_fd_sc_hs__a21o_2
X_5160_ _0630_ _2501_ VSS VSS VCC VCC _2502_ sky130_fd_sc_hs__xnor2_1
X_5091_ _0776_ _2428_ _2293_ VSS VSS VCC VCC _2439_ sky130_fd_sc_hs__o21ai_1
X_4111_ _1728_ VSS VSS VCC VCC _0103_ sky130_fd_sc_hs__clkbuf_1
X_4042_ u_bits.i_op2\[21\] u_bits.i_op2\[19\] _1681_ VSS VSS VCC VCC _1686_
+ sky130_fd_sc_hs__mux2_1
X_4944_ _2064_ _2289_ VSS VSS VCC VCC _2304_ sky130_fd_sc_hs__nor2_1
X_4875_ _2161_ _2269_ u_muldiv.o_div\[29\] VSS VSS VCC VCC _2270_ sky130_fd_sc_hs__a21oi_1
X_3826_ _0784_ _0787_ _0780_ _0795_ _0788_ _0789_ VSS VSS VCC VCC _1546_ sky130_fd_sc_hs__mux4_1
X_3757_ u_muldiv.mul\[12\] _0748_ _1400_ VSS VSS VCC VCC _1482_ sky130_fd_sc_hs__o21ai_1
X_2708_ _0502_ _0507_ _0510_ _0521_ _0522_ VSS VSS VCC VCC _0523_ sky130_fd_sc_hs__o221a_1
X_3688_ _1416_ _1417_ _1336_ u_pc_sel.i_pc_next\[7\] VSS VSS VCC VCC o_result[7]
+ sky130_fd_sc_hs__a2bb2o_2
X_2639_ _0453_ VSS VSS VCC VCC _0454_ sky130_fd_sc_hs__buf_2
X_5427_ clknet_leaf_52_i_clk _0075_ VSS VSS VCC VCC u_bits.i_op2\[18\] sky130_fd_sc_hs__dfxtp_4
X_5358_ clknet_leaf_40_i_clk _0006_ VSS VSS VCC VCC u_muldiv.mul\[54\] sky130_fd_sc_hs__dfxtp_1
X_4309_ _1832_ VSS VSS VCC VCC _1833_ sky130_fd_sc_hs__clkbuf_4
X_5289_ u_muldiv.divisor\[5\] _2284_ _2285_ u_muldiv.divisor\[6\] VSS VSS VCC
+ VCC _0396_ sky130_fd_sc_hs__a22o_1
X_2990_ _0629_ _0769_ _0714_ VSS VSS VCC VCC _0803_ sky130_fd_sc_hs__a21oi_1
X_4660_ _2042_ _2043_ _2081_ _2040_ _2082_ VSS VSS VCC VCC _2083_ sky130_fd_sc_hs__o311a_1
X_3611_ _0998_ _1344_ _0879_ VSS VSS VCC VCC _1345_ sky130_fd_sc_hs__mux2_1
X_4591_ op_cnt\[0\] op_cnt\[1\] _2018_ VSS VSS VCC VCC _0293_ sky130_fd_sc_hs__o21a_1
X_3542_ _1275_ _1276_ _1278_ _0744_ VSS VSS VCC VCC _1279_ sky130_fd_sc_hs__o2bb2a_1
X_3473_ _1227_ VSS VSS VCC VCC o_wdata[18] sky130_fd_sc_hs__buf_2
X_5212_ _0943_ _2362_ _2548_ VSS VSS VCC VCC _2549_ sky130_fd_sc_hs__and3_1
X_5143_ _2486_ VSS VSS VCC VCC _0377_ sky130_fd_sc_hs__clkbuf_1
X_5074_ u_muldiv.dividend\[13\] u_muldiv.dividend\[12\] _2403_ VSS VSS VCC VCC
+ _2423_ sky130_fd_sc_hs__or3_2
X_4025_ u_bits.i_op2\[16\] u_bits.i_op2\[14\] _1657_ VSS VSS VCC VCC _1674_
+ sky130_fd_sc_hs__mux2_1
X_4927_ _1839_ VSS VSS VCC VCC _2288_ sky130_fd_sc_hs__clkbuf_4
X_4858_ _2181_ _2254_ _2256_ VSS VSS VCC VCC _0322_ sky130_fd_sc_hs__a21oi_1
X_3809_ u_bits.i_op2\[16\] _0653_ VSS VSS VCC VCC _1530_ sky130_fd_sc_hs__nand2_1
X_4789_ u_muldiv.o_div\[11\] u_muldiv.o_div\[12\] _2194_ VSS VSS VCC VCC _2201_
+ sky130_fd_sc_hs__or3_2
X_5761_ clknet_leaf_19_i_clk _0404_ VSS VSS VCC VCC u_muldiv.divisor\[13\]
+ sky130_fd_sc_hs__dfxtp_1
X_2973_ u_bits.i_op1\[6\] VSS VSS VCC VCC _0786_ sky130_fd_sc_hs__clkbuf_4
X_4712_ _2030_ _2131_ _2132_ _2133_ _2134_ VSS VSS VCC VCC _2135_ sky130_fd_sc_hs__a311oi_4
X_5692_ clknet_leaf_26_i_clk _0335_ VSS VSS VCC VCC u_muldiv.quotient_msk\[6\]
+ sky130_fd_sc_hs__dfxtp_1
X_4643_ u_muldiv.divisor\[3\] u_muldiv.dividend\[3\] VSS VSS VCC VCC _2066_
+ sky130_fd_sc_hs__and2b_1
X_4574_ _2012_ VSS VSS VCC VCC _0282_ sky130_fd_sc_hs__clkbuf_1
X_3525_ _1261_ _0693_ _0758_ VSS VSS VCC VCC _1262_ sky130_fd_sc_hs__mux2_1
X_3456_ _1218_ VSS VSS VCC VCC o_wdata[10] sky130_fd_sc_hs__buf_2
X_3387_ _0610_ _1164_ _0494_ VSS VSS VCC VCC _1165_ sky130_fd_sc_hs__o21a_2
X_5126_ _2385_ _2469_ _0647_ VSS VSS VCC VCC _2471_ sky130_fd_sc_hs__a21o_1
X_5057_ _2405_ _2406_ _2407_ VSS VSS VCC VCC _2408_ sky130_fd_sc_hs__o21ai_1
X_4008_ u_bits.i_op2\[11\] u_bits.i_op2\[9\] _1657_ VSS VSS VCC VCC _1662_
+ sky130_fd_sc_hs__mux2_1
X_3310_ _1070_ _1094_ _1103_ VSS VSS VCC VCC _1104_ sky130_fd_sc_hs__a21oi_2
X_4290_ csr_data\[27\] i_csr_data[27] _1811_ VSS VSS VCC VCC _1820_ sky130_fd_sc_hs__mux2_1
X_3241_ _0750_ o_add[28] _1039_ VSS VSS VCC VCC _1040_ sky130_fd_sc_hs__a21o_1
X_3172_ _0920_ _0973_ _0974_ VSS VSS VCC VCC _0975_ sky130_fd_sc_hs__a21o_1
X_5744_ clknet_leaf_21_i_clk _0387_ VSS VSS VCC VCC u_muldiv.dividend\[28\]
+ sky130_fd_sc_hs__dfxtp_4
X_2956_ _0768_ u_bits.i_op2\[21\] VSS VSS VCC VCC _0769_ sky130_fd_sc_hs__nand2_1
X_5675_ clknet_leaf_31_i_clk _0318_ VSS VSS VCC VCC u_muldiv.o_div\[21\] sky130_fd_sc_hs__dfxtp_1
X_2887_ u_bits.i_op1\[31\] VSS VSS VCC VCC _0702_ sky130_fd_sc_hs__buf_4
X_4626_ u_muldiv.dividend\[10\] u_muldiv.divisor\[10\] VSS VSS VCC VCC _2049_
+ sky130_fd_sc_hs__or2b_1
X_4557_ _1150_ _2006_ VSS VSS VCC VCC _0271_ sky130_fd_sc_hs__nor2_1
X_4488_ u_muldiv.mul\[4\] u_muldiv.mul\[5\] _1584_ VSS VSS VCC VCC _1975_
+ sky130_fd_sc_hs__mux2_1
X_3508_ _1244_ _1245_ VSS VSS VCC VCC o_wsel[3] sky130_fd_sc_hs__nor2_4
X_3439_ _1206_ VSS VSS VCC VCC _1207_ sky130_fd_sc_hs__buf_4
X_5109_ u_muldiv.dividend\[15\] _2455_ _2378_ VSS VSS VCC VCC _2456_ sky130_fd_sc_hs__mux2_1
X_3790_ _0861_ _0862_ _1339_ _1343_ _0789_ _0674_ VSS VSS VCC VCC _1512_ sky130_fd_sc_hs__mux4_1
X_2810_ _0617_ VSS VSS VCC VCC _0625_ sky130_fd_sc_hs__inv_2
X_2741_ _0554_ _0555_ VSS VSS VCC VCC _0556_ sky130_fd_sc_hs__xnor2_2
X_5460_ clknet_leaf_10_i_clk _0108_ VSS VSS VCC VCC o_pc_target[2] sky130_fd_sc_hs__dfxtp_2
X_2672_ u_bits.i_op1\[17\] u_muldiv.add_prev\[17\] _0450_ VSS VSS VCC VCC
+ _0487_ sky130_fd_sc_hs__mux2_1
X_4411_ _1916_ _1917_ _1833_ VSS VSS VCC VCC _1918_ sky130_fd_sc_hs__a21oi_1
X_5391_ clknet_leaf_49_i_clk _0039_ VSS VSS VCC VCC u_bits.i_op1\[23\] sky130_fd_sc_hs__dfxtp_2
X_4342_ _1860_ _1861_ VSS VSS VCC VCC _1862_ sky130_fd_sc_hs__nor2_1
X_4273_ _1711_ VSS VSS VCC VCC _1811_ sky130_fd_sc_hs__clkbuf_4
X_3224_ _1017_ _1023_ VSS VSS VCC VCC _1024_ sky130_fd_sc_hs__xnor2_2


