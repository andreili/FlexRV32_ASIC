* NGSPICE file created from rv_ctrl.ext - technology: sky130A

X_66_ o_decode_stall VSS VSS VCC VCC o_fetch_stall sky130_fd_sc_hs__buf_2
X_49_ _12_ _19_ _21_ VSS VSS VCC VCC _22_ sky130_fd_sc_hs__a21o_1
X_65_ o_alu2_flush VSS VSS VCC VCC o_decode_flush sky130_fd_sc_hs__buf_2
X_48_ i_alu1_rd[2] _20_ i_alu1_mem_rd VSS VSS VCC VCC _21_ sky130_fd_sc_hs__o21ai_1
X_64_ clknet_1_0__leaf_i_clk _01_ VSS VSS VCC VCC inst_sup\[1\] sky130_fd_sc_hs__dfxtp_1
X_47_ i_alu1_rd[1] i_alu1_rd[0] i_alu1_rd[3] i_alu1_rd[4] VSS VSS VCC VCC
+ _20_ sky130_fd_sc_hs__or4_1
X_63_ clknet_1_1__leaf_i_clk _00_ VSS VSS VCC VCC inst_sup\[0\] sky130_fd_sc_hs__dfxtp_1
X_46_ _13_ _16_ _17_ _18_ VSS VSS VCC VCC _19_ sky130_fd_sc_hs__or4b_1
X_29_ i_decode_rs1[2] VSS VSS VCC VCC _02_ sky130_fd_sc_hs__inv_2
X_62_ inst_sup\[1\] o_decode_stall _28_ VSS VSS VCC VCC _01_ sky130_fd_sc_hs__a21o_1
X_45_ _04_ i_decode_rs2[1] _14_ i_alu1_rd[2] VSS VSS VCC VCC _18_ sky130_fd_sc_hs__o22a_1
Xclkbuf_0_i_clk i_clk VSS VSS VCC VCC clknet_0_i_clk sky130_fd_sc_hs__clkbuf_16
X_61_ inst_sup\[0\] i_alu2_ready _22_ _23_ o_alu2_flush VSS VSS VCC VCC _28_
+ sky130_fd_sc_hs__a41o_1
X_44_ i_alu1_rd[3] i_decode_rs2[3] VSS VSS VCC VCC _17_ sky130_fd_sc_hs__xor2_1
X_60_ inst_sup\[0\] o_decode_stall _27_ VSS VSS VCC VCC _00_ sky130_fd_sc_hs__a21o_1
X_43_ _04_ i_decode_rs2[1] _14_ i_alu1_rd[2] _15_ VSS VSS VCC VCC _16_ sky130_fd_sc_hs__a221o_1
X_42_ i_alu1_rd[4] i_decode_rs2[4] VSS VSS VCC VCC _15_ sky130_fd_sc_hs__xor2_1
X_41_ i_decode_rs2[2] VSS VSS VCC VCC _14_ sky130_fd_sc_hs__inv_2
X_40_ i_alu1_rd[0] i_decode_rs2[0] VSS VSS VCC VCC _13_ sky130_fd_sc_hs__xor2_1
X_59_ i_decode_inst_sup i_alu2_ready _22_ _23_ o_alu2_flush VSS VSS VCC VCC
+ _27_ sky130_fd_sc_hs__a41o_1
X_58_ _26_ VSS VSS VCC VCC o_alu1_flush sky130_fd_sc_hs__buf_2
X_57_ o_alu2_flush _25_ VSS VSS VCC VCC _26_ sky130_fd_sc_hs__or2_1
X_56_ _22_ _23_ o_alu1_stall VSS VSS VCC VCC _25_ sky130_fd_sc_hs__a21oi_1
X_39_ _03_ _05_ _09_ _11_ VSS VSS VCC VCC _12_ sky130_fd_sc_hs__or4b_1
X_55_ _24_ VSS VSS VCC VCC o_alu2_flush sky130_fd_sc_hs__clkbuf_4
X_38_ _06_ i_decode_rs1[3] i_decode_rs1[4] _07_ _10_ VSS VSS VCC VCC _11_
+ sky130_fd_sc_hs__o221a_1
X_54_ i_pc_change i_reset_n VSS VSS VCC VCC _24_ sky130_fd_sc_hs__or2b_1
X_37_ i_decode_rs1[1] i_alu1_rd[1] VSS VSS VCC VCC _10_ sky130_fd_sc_hs__or2b_1
X_53_ inst_sup\[1\] VSS VSS VCC VCC o_inv_inst sky130_fd_sc_hs__inv_2
X_36_ _06_ i_decode_rs1[3] i_decode_rs1[4] _07_ _08_ VSS VSS VCC VCC _09_
+ sky130_fd_sc_hs__a221o_1
Xclkbuf_1_1__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_1_1__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_52_ i_alu2_ready VSS VSS VCC VCC o_alu1_stall sky130_fd_sc_hs__inv_2
X_35_ i_alu1_rd[0] i_decode_rs1[0] VSS VSS VCC VCC _08_ sky130_fd_sc_hs__xor2_1
X_51_ i_alu2_ready _22_ _23_ VSS VSS VCC VCC o_decode_stall sky130_fd_sc_hs__nand3_4
X_34_ i_alu1_rd[4] VSS VSS VCC VCC _07_ sky130_fd_sc_hs__inv_2
X_50_ i_need_pause i_reset_n VSS VSS VCC VCC _23_ sky130_fd_sc_hs__nor2b_2
X_33_ i_alu1_rd[3] VSS VSS VCC VCC _06_ sky130_fd_sc_hs__inv_2
X_32_ _04_ i_decode_rs1[1] _02_ i_alu1_rd[2] VSS VSS VCC VCC _05_ sky130_fd_sc_hs__a22o_1
X_31_ i_alu1_rd[1] VSS VSS VCC VCC _04_ sky130_fd_sc_hs__inv_2
X_30_ i_alu1_rd[2] _02_ VSS VSS VCC VCC _03_ sky130_fd_sc_hs__nor2_1
Xclkbuf_1_0__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_1_0__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16

