* NGSPICE file created from rv_fetch.ext - technology: sky130A

X_0985_ _0059_ VSS VSS VCC VCC _0029_ sky130_fd_sc_hs__clkbuf_1
X_0419_ _0072_ VSS VSS VCC VCC o_instruction[19] sky130_fd_sc_hs__buf_2
X_0770_ o_pc[5] _0287_ VSS VSS VCC VCC _0295_ sky130_fd_sc_hs__and2_1
X_0968_ u_buf.data\[0\]\[21\] u_buf.latch_hi\[5\] _0045_ VSS VSS VCC VCC _0051_
+ sky130_fd_sc_hs__mux2_1
X_0899_ u_buf.is_head\[4\] _0378_ _0379_ u_buf.is_head\[2\] VSS VSS VCC VCC
+ _0381_ sky130_fd_sc_hs__a22o_1
X_0822_ _0264_ _0339_ _0340_ VSS VSS VCC VCC _0341_ sky130_fd_sc_hs__and3_1
X_0684_ i_instruction[15] _0223_ _0224_ u_buf.data\[0\]\[15\] VSS VSS VCC VCC
+ _0230_ sky130_fd_sc_hs__a22o_1
X_0753_ o_pc[2] _0267_ o_pc[3] VSS VSS VCC VCC _0280_ sky130_fd_sc_hs__a21o_1
X_1167_ clknet_4_10_0_i_clk o_pc_next[11] VSS VSS VCC VCC o_pc[11] sky130_fd_sc_hs__dfxtp_4
X_1098_ clknet_4_0_0_i_clk u_buf.g_data\[0\].d_next\[5\] VSS VSS VCC VCC u_buf.data\[0\]\[5\]
+ sky130_fd_sc_hs__dfxtp_1
X_1021_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[27\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[27\] sky130_fd_sc_hs__dfxtp_1
X_0805_ o_pc[5] _0287_ _0324_ o_pc[9] VSS VSS VCC VCC _0326_ sky130_fd_sc_hs__a31o_1
X_0736_ _0106_ VSS VSS VCC VCC _0265_ sky130_fd_sc_hs__inv_2
X_0667_ i_instruction[8] _0209_ _0211_ u_buf.data\[0\]\[8\] VSS VSS VCC VCC
+ _0220_ sky130_fd_sc_hs__a22o_1
X_0598_ u_buf.data\[1\]\[11\] _0178_ _0175_ i_instruction[11] _0179_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[11\] sky130_fd_sc_hs__a221o_1
X_0521_ u_buf.data\[3\]\[13\] _0129_ _0123_ VSS VSS VCC VCC _0133_ sky130_fd_sc_hs__and3_1
X_0452_ u_buf.data\[0\]\[3\] u_buf.latch_hi\[3\] _0088_ VSS VSS VCC VCC _0090_
+ sky130_fd_sc_hs__mux2_1
X_1004_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[10\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[10\] sky130_fd_sc_hs__dfxtp_1
X_0719_ i_instruction[31] _0206_ _0210_ u_buf.data\[0\]\[31\] VSS VSS VCC VCC
+ _0249_ sky130_fd_sc_hs__a22o_1
X_0435_ u_buf.data\[0\]\[27\] u_buf.data\[0\]\[11\] _0077_ VSS VSS VCC VCC
+ _0081_ sky130_fd_sc_hs__mux2_1
X_0504_ u_buf.data\[2\]\[6\] _0109_ _0112_ i_instruction[6] _0122_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[6\] sky130_fd_sc_hs__a221o_1
X_0984_ u_buf.data\[0\]\[29\] u_buf.latch_hi\[13\] _0250_ VSS VSS VCC VCC
+ _0059_ sky130_fd_sc_hs__mux2_1
X_0418_ u_buf.data\[0\]\[19\] u_buf.data\[0\]\[3\] _0068_ VSS VSS VCC VCC
+ _0072_ sky130_fd_sc_hs__mux2_1
X_0967_ _0050_ VSS VSS VCC VCC _0020_ sky130_fd_sc_hs__clkbuf_1
X_0898_ _0378_ _0379_ VSS VSS VCC VCC _0380_ sky130_fd_sc_hs__nor2_1
X_0752_ o_pc[2] o_pc[3] _0267_ VSS VSS VCC VCC _0279_ sky130_fd_sc_hs__nand3_1
X_0821_ o_pc[10] o_pc[11] _0325_ VSS VSS VCC VCC _0340_ sky130_fd_sc_hs__nand3_1
X_0683_ u_buf.data\[1\]\[14\] _0222_ _0229_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[14\]
+ sky130_fd_sc_hs__a21o_1
X_1166_ clknet_4_10_0_i_clk o_pc_next[10] VSS VSS VCC VCC o_pc[10] sky130_fd_sc_hs__dfxtp_4
X_1097_ clknet_4_0_0_i_clk u_buf.g_data\[0\].d_next\[4\] VSS VSS VCC VCC u_buf.data\[0\]\[4\]
+ sky130_fd_sc_hs__dfxtp_1
X_1020_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[26\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[26\] sky130_fd_sc_hs__dfxtp_1
X_0735_ _0263_ VSS VSS VCC VCC _0264_ sky130_fd_sc_hs__buf_2
X_0804_ o_pc[5] o_pc[9] _0287_ _0324_ VSS VSS VCC VCC _0325_ sky130_fd_sc_hs__and4_1
X_0666_ u_buf.data\[1\]\[7\] _0208_ _0219_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[7\]
+ sky130_fd_sc_hs__a21o_1
X_0597_ u_buf.data\[2\]\[11\] _0173_ _0176_ VSS VSS VCC VCC _0179_ sky130_fd_sc_hs__and3_1
X_1149_ clknet_4_2_0_i_clk _0025_ VSS VSS VCC VCC u_buf.latch_hi\[9\] sky130_fd_sc_hs__dfxtp_1
X_0520_ u_buf.data\[2\]\[12\] _0127_ _0128_ i_instruction[12] _0132_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[12\] sky130_fd_sc_hs__a221o_1
X_0451_ _0089_ VSS VSS VCC VCC o_instruction[2] sky130_fd_sc_hs__buf_2
X_1003_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[9\] VSS VSS VCC VCC u_buf.data\[3\]\[9\]
+ sky130_fd_sc_hs__dfxtp_1
X_0718_ u_buf.data\[1\]\[30\] _0207_ _0248_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[30\]
+ sky130_fd_sc_hs__a21o_1
X_0649_ _0107_ _0205_ VSS VSS VCC VCC _0210_ sky130_fd_sc_hs__nor2_2
Xclkbuf_4_15_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_15_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0434_ _0080_ VSS VSS VCC VCC o_instruction[26] sky130_fd_sc_hs__buf_2
X_0503_ u_buf.data\[3\]\[6\] _0113_ _0115_ VSS VSS VCC VCC _0122_ sky130_fd_sc_hs__and3_1
X_0983_ _0058_ VSS VSS VCC VCC _0028_ sky130_fd_sc_hs__clkbuf_1
X_0417_ _0071_ VSS VSS VCC VCC o_instruction[18] sky130_fd_sc_hs__buf_2
X_0966_ u_buf.data\[0\]\[20\] u_buf.latch_hi\[4\] _0045_ VSS VSS VCC VCC _0050_
+ sky130_fd_sc_hs__mux2_1
X_0897_ u_buf.i_push _0204_ VSS VSS VCC VCC _0379_ sky130_fd_sc_hs__and2_1
X_0751_ _0255_ i_pc_trap[3] _0277_ _0065_ VSS VSS VCC VCC _0278_ sky130_fd_sc_hs__o211a_1
X_0820_ o_pc[10] _0325_ o_pc[11] VSS VSS VCC VCC _0339_ sky130_fd_sc_hs__a21o_1
X_0682_ i_instruction[14] _0223_ _0224_ u_buf.data\[0\]\[14\] VSS VSS VCC VCC
+ _0229_ sky130_fd_sc_hs__a22o_1
X_1165_ clknet_4_10_0_i_clk o_pc_next[9] VSS VSS VCC VCC o_pc[9] sky130_fd_sc_hs__dfxtp_4
X_1096_ clknet_4_0_0_i_clk u_buf.g_data\[0\].d_next\[3\] VSS VSS VCC VCC u_buf.data\[0\]\[3\]
+ sky130_fd_sc_hs__dfxtp_1
X_0949_ _0039_ VSS VSS VCC VCC _0013_ sky130_fd_sc_hs__clkbuf_1
X_0734_ u_buf.first_half _0251_ _0262_ VSS VSS VCC VCC _0263_ sky130_fd_sc_hs__and3b_1
X_0803_ o_pc[6] o_pc[7] o_pc[8] VSS VSS VCC VCC _0324_ sky130_fd_sc_hs__and3_1
X_0665_ i_instruction[7] _0209_ _0211_ u_buf.data\[0\]\[7\] VSS VSS VCC VCC
+ _0219_ sky130_fd_sc_hs__a22o_1
X_0596_ _0158_ VSS VSS VCC VCC _0178_ sky130_fd_sc_hs__buf_2
X_1148_ clknet_4_0_0_i_clk _0024_ VSS VSS VCC VCC u_buf.latch_hi\[8\] sky130_fd_sc_hs__dfxtp_1
X_1079_ clknet_4_12_0_i_clk u_buf.g_data\[1\].d_next\[19\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[19\] sky130_fd_sc_hs__dfxtp_1
X_0450_ u_buf.data\[0\]\[2\] u_buf.latch_hi\[2\] _0088_ VSS VSS VCC VCC _0089_
+ sky130_fd_sc_hs__mux2_1
Xclkbuf_4_11_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_11_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_1002_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[8\] VSS VSS VCC VCC u_buf.data\[3\]\[8\]
+ sky130_fd_sc_hs__dfxtp_1
X_0648_ _0206_ VSS VSS VCC VCC _0209_ sky130_fd_sc_hs__buf_2
X_0717_ i_instruction[30] _0206_ _0210_ u_buf.data\[0\]\[30\] VSS VSS VCC VCC
+ _0248_ sky130_fd_sc_hs__a22o_1
X_0579_ u_buf.data\[2\]\[4\] _0161_ _0162_ VSS VSS VCC VCC _0168_ sky130_fd_sc_hs__and3_1
X_0502_ u_buf.data\[2\]\[5\] _0109_ _0112_ i_instruction[5] _0121_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[5\] sky130_fd_sc_hs__a221o_1
X_0433_ u_buf.data\[0\]\[26\] u_buf.data\[0\]\[10\] _0077_ VSS VSS VCC VCC
+ _0080_ sky130_fd_sc_hs__mux2_1
X_0982_ u_buf.data\[0\]\[28\] u_buf.latch_hi\[12\] _0250_ VSS VSS VCC VCC
+ _0058_ sky130_fd_sc_hs__mux2_1
X_0416_ u_buf.data\[0\]\[18\] u_buf.data\[0\]\[2\] _0068_ VSS VSS VCC VCC
+ _0071_ sky130_fd_sc_hs__mux2_1
X_0965_ _0049_ VSS VSS VCC VCC _0019_ sky130_fd_sc_hs__clkbuf_1
X_0896_ u_buf.i_push _0204_ VSS VSS VCC VCC _0378_ sky130_fd_sc_hs__nor2_1
X_0750_ _0270_ i_pc_target[3] _0275_ _0276_ i_ebreak VSS VSS VCC VCC _0277_
+ sky130_fd_sc_hs__a221o_1
X_0681_ u_buf.data\[1\]\[13\] _0222_ _0228_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[13\]
+ sky130_fd_sc_hs__a21o_1
X_1164_ clknet_4_10_0_i_clk o_pc_next[8] VSS VSS VCC VCC o_pc[8] sky130_fd_sc_hs__dfxtp_4
X_1095_ clknet_4_0_0_i_clk u_buf.g_data\[0\].d_next\[2\] VSS VSS VCC VCC u_buf.data\[0\]\[2\]
+ sky130_fd_sc_hs__dfxtp_1
X_0948_ o_addr[13] _0354_ _0395_ VSS VSS VCC VCC _0039_ sky130_fd_sc_hs__mux2_1
X_0879_ u_buf.data\[3\]\[18\] _0373_ _0374_ i_instruction[18] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[18\] sky130_fd_sc_hs__a22o_1
X_0802_ _0254_ i_pc_trap[9] _0321_ _0322_ i_reset_n VSS VSS VCC VCC _0323_
+ sky130_fd_sc_hs__o221a_1
X_0733_ _0250_ VSS VSS VCC VCC _0262_ sky130_fd_sc_hs__inv_2
X_0664_ u_buf.data\[1\]\[6\] _0208_ _0218_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[6\]
+ sky130_fd_sc_hs__a21o_1
X_0595_ u_buf.data\[1\]\[10\] _0164_ _0175_ i_instruction[10] _0177_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[10\] sky130_fd_sc_hs__a221o_1
X_1078_ clknet_4_5_0_i_clk u_buf.g_data\[1\].d_next\[18\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[18\] sky130_fd_sc_hs__dfxtp_1
X_1147_ clknet_4_0_0_i_clk _0023_ VSS VSS VCC VCC u_buf.latch_hi\[7\] sky130_fd_sc_hs__dfxtp_1
X_1001_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[7\] VSS VSS VCC VCC u_buf.data\[3\]\[7\]
+ sky130_fd_sc_hs__dfxtp_1
X_0578_ u_buf.data\[1\]\[3\] _0164_ _0160_ i_instruction[3] _0167_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[3\] sky130_fd_sc_hs__a221o_1
X_0647_ _0207_ VSS VSS VCC VCC _0208_ sky130_fd_sc_hs__buf_2
X_0716_ u_buf.data\[1\]\[29\] _0235_ _0247_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[29\]
+ sky130_fd_sc_hs__a21o_1
X_0432_ _0079_ VSS VSS VCC VCC o_instruction[25] sky130_fd_sc_hs__buf_2
X_0501_ u_buf.data\[3\]\[5\] _0113_ _0115_ VSS VSS VCC VCC _0121_ sky130_fd_sc_hs__and3_1
Xclkbuf_4_9_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_9_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0981_ _0057_ VSS VSS VCC VCC _0027_ sky130_fd_sc_hs__clkbuf_1
X_0415_ _0070_ VSS VSS VCC VCC o_instruction[17] sky130_fd_sc_hs__buf_2
X_0964_ u_buf.data\[0\]\[19\] u_buf.latch_hi\[3\] _0045_ VSS VSS VCC VCC _0049_
+ sky130_fd_sc_hs__mux2_1
X_0895_ i_reset_n _0063_ VSS VSS VCC VCC _0377_ sky130_fd_sc_hs__nand2_2
X_0680_ i_instruction[13] _0223_ _0224_ u_buf.data\[0\]\[13\] VSS VSS VCC VCC
+ _0228_ sky130_fd_sc_hs__a22o_1
X_1163_ clknet_4_10_0_i_clk o_pc_next[7] VSS VSS VCC VCC o_pc[7] sky130_fd_sc_hs__dfxtp_4
X_1094_ clknet_4_3_0_i_clk u_buf.g_data\[0\].d_next\[1\] VSS VSS VCC VCC u_buf.data\[0\]\[1\]
+ sky130_fd_sc_hs__dfxtp_1
X_0947_ o_addr[12] _0391_ _0037_ _0038_ VSS VSS VCC VCC _0012_ sky130_fd_sc_hs__a22o_1
X_0878_ u_buf.data\[3\]\[17\] _0373_ _0374_ i_instruction[17] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[17\] sky130_fd_sc_hs__a22o_1
X_0801_ _0270_ i_pc_target[9] _0258_ VSS VSS VCC VCC _0322_ sky130_fd_sc_hs__a21o_1
X_0732_ u_buf.data\[0\]\[0\] u_buf.data\[0\]\[1\] VSS VSS VCC VCC _0261_ sky130_fd_sc_hs__nand2_1
X_0663_ i_instruction[6] _0209_ _0211_ u_buf.data\[0\]\[6\] VSS VSS VCC VCC
+ _0218_ sky130_fd_sc_hs__a22o_1
X_0594_ u_buf.data\[2\]\[10\] _0173_ _0176_ VSS VSS VCC VCC _0177_ sky130_fd_sc_hs__and3_1
X_1146_ clknet_4_0_0_i_clk _0022_ VSS VSS VCC VCC u_buf.latch_hi\[6\] sky130_fd_sc_hs__dfxtp_1
X_1077_ clknet_4_13_0_i_clk u_buf.g_data\[1\].d_next\[17\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[17\] sky130_fd_sc_hs__dfxtp_1
X_1000_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[6\] VSS VSS VCC VCC u_buf.data\[3\]\[6\]
+ sky130_fd_sc_hs__dfxtp_1
X_0715_ i_instruction[29] _0236_ _0237_ u_buf.data\[0\]\[29\] VSS VSS VCC VCC
+ _0247_ sky130_fd_sc_hs__a22o_1
X_0646_ _0204_ _0206_ VSS VSS VCC VCC _0207_ sky130_fd_sc_hs__nor2_1
X_0577_ u_buf.data\[2\]\[3\] _0161_ _0162_ VSS VSS VCC VCC _0167_ sky130_fd_sc_hs__and3_1
Xclkbuf_4_5_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_5_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_1129_ clknet_4_11_0_i_clk _0005_ VSS VSS VCC VCC o_addr[5] sky130_fd_sc_hs__dfxtp_2
X_0431_ u_buf.data\[0\]\[25\] u_buf.data\[0\]\[9\] _0077_ VSS VSS VCC VCC
+ _0079_ sky130_fd_sc_hs__mux2_1
X_0500_ u_buf.data\[2\]\[4\] _0109_ _0112_ i_instruction[4] _0120_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[4\] sky130_fd_sc_hs__a221o_1
X_0629_ u_buf.data\[2\]\[25\] _0187_ _0190_ VSS VSS VCC VCC _0197_ sky130_fd_sc_hs__and3_1
Xclkbuf_0_i_clk i_clk VSS VSS VCC VCC clknet_0_i_clk sky130_fd_sc_hs__clkbuf_16
X_0980_ u_buf.data\[0\]\[27\] u_buf.latch_hi\[11\] _0250_ VSS VSS VCC VCC
+ _0057_ sky130_fd_sc_hs__mux2_1
X_0414_ u_buf.data\[0\]\[17\] u_buf.data\[0\]\[1\] _0068_ VSS VSS VCC VCC
+ _0070_ sky130_fd_sc_hs__mux2_1
X_0963_ _0048_ VSS VSS VCC VCC _0018_ sky130_fd_sc_hs__clkbuf_1
X_0894_ u_buf.data\[3\]\[31\] _0369_ _0371_ i_instruction[31] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[31\] sky130_fd_sc_hs__a22o_1
X_1162_ clknet_4_10_0_i_clk o_pc_next[6] VSS VSS VCC VCC o_pc[6] sky130_fd_sc_hs__dfxtp_4
X_1093_ clknet_4_2_0_i_clk u_buf.g_data\[0\].d_next\[0\] VSS VSS VCC VCC u_buf.data\[0\]\[0\]
+ sky130_fd_sc_hs__dfxtp_1
X_0877_ u_buf.data\[3\]\[16\] _0373_ _0374_ i_instruction[16] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[16\] sky130_fd_sc_hs__a22o_1
X_0946_ _0346_ _0391_ VSS VSS VCC VCC _0038_ sky130_fd_sc_hs__nor2_1
X_0731_ _0255_ i_pc_trap[1] _0259_ _0065_ VSS VSS VCC VCC _0260_ sky130_fd_sc_hs__o211a_1
X_0800_ _0270_ _0319_ _0320_ VSS VSS VCC VCC _0321_ sky130_fd_sc_hs__nor3b_1
X_0662_ u_buf.data\[1\]\[5\] _0208_ _0217_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[5\]
+ sky130_fd_sc_hs__a21o_1
X_0593_ _0157_ VSS VSS VCC VCC _0176_ sky130_fd_sc_hs__clkbuf_2
X_1145_ clknet_4_0_0_i_clk _0021_ VSS VSS VCC VCC u_buf.latch_hi\[5\] sky130_fd_sc_hs__dfxtp_1
X_1076_ clknet_4_5_0_i_clk u_buf.g_data\[1\].d_next\[16\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[16\] sky130_fd_sc_hs__dfxtp_1
Xclkbuf_4_1_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_1_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0929_ o_addr[6] _0301_ _0395_ VSS VSS VCC VCC _0398_ sky130_fd_sc_hs__mux2_1
X_0645_ u_buf.is_head\[1\] _0107_ _0205_ VSS VSS VCC VCC _0206_ sky130_fd_sc_hs__a21o_1
X_0714_ u_buf.data\[1\]\[28\] _0235_ _0246_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[28\]
+ sky130_fd_sc_hs__a21o_1
X_0576_ u_buf.data\[1\]\[2\] _0164_ _0160_ i_instruction[2] _0166_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[2\] sky130_fd_sc_hs__a221o_1
X_1128_ clknet_4_8_0_i_clk _0004_ VSS VSS VCC VCC o_addr[4] sky130_fd_sc_hs__dfxtp_4
X_1059_ clknet_4_11_0_i_clk u_buf.g_data\[1\].h_next VSS VSS VCC VCC u_buf.is_head\[2\]
+ sky130_fd_sc_hs__dfxtp_1
X_0430_ _0078_ VSS VSS VCC VCC o_instruction[24] sky130_fd_sc_hs__buf_2
X_0628_ u_buf.data\[1\]\[24\] _0192_ _0189_ i_instruction[24] _0196_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[24\] sky130_fd_sc_hs__a221o_1
X_0559_ u_buf.data\[3\]\[30\] _0110_ _0114_ VSS VSS VCC VCC _0154_ sky130_fd_sc_hs__and3_1
X_0413_ _0069_ VSS VSS VCC VCC o_instruction[16] sky130_fd_sc_hs__buf_2
X_0962_ u_buf.data\[0\]\[18\] u_buf.latch_hi\[2\] _0045_ VSS VSS VCC VCC _0048_
+ sky130_fd_sc_hs__mux2_1
X_0893_ u_buf.data\[3\]\[30\] _0369_ _0371_ i_instruction[30] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[30\] sky130_fd_sc_hs__a22o_1
X_1161_ clknet_4_10_0_i_clk o_pc_next[5] VSS VSS VCC VCC o_pc[5] sky130_fd_sc_hs__dfxtp_4
X_1092_ clknet_4_9_0_i_clk u_buf.g_data\[0\].h_next VSS VSS VCC VCC u_buf.is_head\[1\]
+ sky130_fd_sc_hs__dfxtp_1
X_0876_ u_buf.data\[3\]\[15\] _0373_ _0374_ i_instruction[15] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[15\] sky130_fd_sc_hs__a22o_1
X_0945_ _0257_ _0036_ _0347_ VSS VSS VCC VCC _0037_ sky130_fd_sc_hs__o21ai_1
X_0730_ _0257_ i_pc_target[1] _0258_ VSS VSS VCC VCC _0259_ sky130_fd_sc_hs__a21o_1
X_0661_ i_instruction[5] _0209_ _0211_ u_buf.data\[0\]\[5\] VSS VSS VCC VCC
+ _0217_ sky130_fd_sc_hs__a22o_1
X_0592_ _0159_ VSS VSS VCC VCC _0175_ sky130_fd_sc_hs__buf_2
X_1075_ clknet_4_7_0_i_clk u_buf.g_data\[1\].d_next\[15\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[15\] sky130_fd_sc_hs__dfxtp_1
X_1144_ clknet_4_0_0_i_clk _0020_ VSS VSS VCC VCC u_buf.latch_hi\[4\] sky130_fd_sc_hs__dfxtp_1
X_0928_ _0397_ VSS VSS VCC VCC _0005_ sky130_fd_sc_hs__clkbuf_1
X_0859_ u_buf.data\[3\]\[0\] _0370_ _0372_ i_instruction[0] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[0\] sky130_fd_sc_hs__a22o_1
X_0644_ u_buf.i_push u_buf.is_head\[0\] VSS VSS VCC VCC _0205_ sky130_fd_sc_hs__and2_1
X_0713_ i_instruction[28] _0236_ _0237_ u_buf.data\[0\]\[28\] VSS VSS VCC VCC
+ _0246_ sky130_fd_sc_hs__a22o_1
X_0575_ u_buf.data\[2\]\[2\] _0161_ _0162_ VSS VSS VCC VCC _0166_ sky130_fd_sc_hs__and3_1
X_1127_ clknet_4_8_0_i_clk _0003_ VSS VSS VCC VCC o_addr[3] sky130_fd_sc_hs__dfxtp_4
X_1058_ clknet_4_6_0_i_clk u_buf.g_data\[2\].d_next\[31\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[31\] sky130_fd_sc_hs__dfxtp_1
X_0558_ u_buf.data\[2\]\[29\] _0141_ _0142_ i_instruction[29] _0153_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[29\] sky130_fd_sc_hs__a221o_1
X_0627_ u_buf.data\[2\]\[24\] _0187_ _0190_ VSS VSS VCC VCC _0196_ sky130_fd_sc_hs__and3_1
X_0489_ _0107_ VSS VSS VCC VCC _0114_ sky130_fd_sc_hs__buf_2
X_0412_ u_buf.data\[0\]\[16\] u_buf.data\[0\]\[0\] _0068_ VSS VSS VCC VCC
+ _0069_ sky130_fd_sc_hs__mux2_1
X_0961_ _0047_ VSS VSS VCC VCC _0017_ sky130_fd_sc_hs__clkbuf_1
X_0892_ u_buf.data\[3\]\[29\] _0375_ _0376_ i_instruction[29] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[29\] sky130_fd_sc_hs__a22o_1
X_1160_ clknet_4_10_0_i_clk o_pc_next[4] VSS VSS VCC VCC o_pc[4] sky130_fd_sc_hs__dfxtp_4
X_1091_ clknet_4_9_0_i_clk u_buf.g_data\[1\].d_next\[31\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[31\] sky130_fd_sc_hs__dfxtp_1
X_0944_ o_addr[12] _0335_ _0349_ _0319_ VSS VSS VCC VCC _0036_ sky130_fd_sc_hs__a2bb2o_1
X_0875_ u_buf.data\[3\]\[14\] _0373_ _0374_ i_instruction[14] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[14\] sky130_fd_sc_hs__a22o_1
X_0660_ u_buf.data\[1\]\[4\] _0208_ _0216_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[4\]
+ sky130_fd_sc_hs__a21o_1
X_0591_ u_buf.data\[1\]\[9\] _0164_ _0160_ i_instruction[9] _0174_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[9\] sky130_fd_sc_hs__a221o_1
X_1143_ clknet_4_0_0_i_clk _0019_ VSS VSS VCC VCC u_buf.latch_hi\[3\] sky130_fd_sc_hs__dfxtp_1
X_1074_ clknet_4_7_0_i_clk u_buf.g_data\[1\].d_next\[14\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[14\] sky130_fd_sc_hs__dfxtp_1
X_0927_ o_addr[5] _0294_ _0395_ VSS VSS VCC VCC _0397_ sky130_fd_sc_hs__mux2_1
X_0789_ _0310_ _0311_ VSS VSS VCC VCC _0312_ sky130_fd_sc_hs__nor2_1
X_0858_ _0371_ VSS VSS VCC VCC _0372_ sky130_fd_sc_hs__buf_2
X_0643_ u_buf.hi_valid _0106_ _0103_ VSS VSS VCC VCC _0204_ sky130_fd_sc_hs__a21o_1
X_0574_ u_buf.data\[1\]\[1\] _0164_ _0160_ i_instruction[1] _0165_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[1\] sky130_fd_sc_hs__a221o_1
X_0712_ u_buf.data\[1\]\[27\] _0235_ _0245_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[27\]
+ sky130_fd_sc_hs__a21o_1
X_1126_ clknet_4_8_0_i_clk _0002_ VSS VSS VCC VCC o_addr[2] sky130_fd_sc_hs__dfxtp_4
X_1057_ clknet_4_12_0_i_clk u_buf.g_data\[2\].d_next\[30\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[30\] sky130_fd_sc_hs__dfxtp_1
X_0557_ u_buf.data\[3\]\[29\] _0143_ _0114_ VSS VSS VCC VCC _0153_ sky130_fd_sc_hs__and3_1
X_0626_ u_buf.data\[1\]\[23\] _0192_ _0189_ i_instruction[23] _0195_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[23\] sky130_fd_sc_hs__a221o_1
X_0488_ _0110_ VSS VSS VCC VCC _0113_ sky130_fd_sc_hs__clkbuf_2
X_1109_ clknet_4_5_0_i_clk u_buf.g_data\[0\].d_next\[16\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[16\] sky130_fd_sc_hs__dfxtp_1
X_0411_ _0067_ VSS VSS VCC VCC _0068_ sky130_fd_sc_hs__clkbuf_4
X_0609_ u_buf.data\[2\]\[17\] _0173_ _0176_ VSS VSS VCC VCC _0185_ sky130_fd_sc_hs__and3_1
X_0960_ u_buf.data\[0\]\[17\] u_buf.latch_hi\[1\] _0045_ VSS VSS VCC VCC _0047_
+ sky130_fd_sc_hs__mux2_1
X_0891_ u_buf.data\[3\]\[28\] _0375_ _0376_ i_instruction[28] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[28\] sky130_fd_sc_hs__a22o_1
X_1090_ clknet_4_12_0_i_clk u_buf.g_data\[1\].d_next\[30\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[30\] sky130_fd_sc_hs__dfxtp_1
X_0874_ u_buf.data\[3\]\[13\] _0373_ _0374_ i_instruction[13] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[13\] sky130_fd_sc_hs__a22o_1
X_0943_ _0035_ VSS VSS VCC VCC _0011_ sky130_fd_sc_hs__clkbuf_1
X_0590_ u_buf.data\[2\]\[9\] _0173_ _0162_ VSS VSS VCC VCC _0174_ sky130_fd_sc_hs__and3_1
X_1142_ clknet_4_0_0_i_clk _0018_ VSS VSS VCC VCC u_buf.latch_hi\[2\] sky130_fd_sc_hs__dfxtp_1
X_1073_ clknet_4_7_0_i_clk u_buf.g_data\[1\].d_next\[13\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[13\] sky130_fd_sc_hs__dfxtp_1
X_0926_ _0396_ VSS VSS VCC VCC _0004_ sky130_fd_sc_hs__clkbuf_1
X_0857_ u_buf.is_head\[4\] _0114_ _0368_ VSS VSS VCC VCC _0371_ sky130_fd_sc_hs__a21o_1
X_0788_ o_pc[7] _0302_ _0264_ VSS VSS VCC VCC _0311_ sky130_fd_sc_hs__o21ai_1
X_0711_ i_instruction[27] _0236_ _0237_ u_buf.data\[0\]\[27\] VSS VSS VCC VCC
+ _0245_ sky130_fd_sc_hs__a22o_1
X_0573_ u_buf.data\[2\]\[1\] _0161_ _0162_ VSS VSS VCC VCC _0165_ sky130_fd_sc_hs__and3_1
X_0642_ u_buf.data\[1\]\[31\] _0158_ _0159_ i_instruction[31] _0203_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[31\] sky130_fd_sc_hs__a221o_1
X_1125_ clknet_4_14_0_i_clk _0001_ VSS VSS VCC VCC o_addr[1] sky130_fd_sc_hs__dfxtp_2
X_1056_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[29\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[29\] sky130_fd_sc_hs__dfxtp_1
X_0909_ u_buf.hi_valid u_buf.is_head\[0\] _0068_ VSS VSS VCC VCC _0387_ sky130_fd_sc_hs__and3b_1
X_0625_ u_buf.data\[2\]\[23\] _0187_ _0190_ VSS VSS VCC VCC _0195_ sky130_fd_sc_hs__and3_1
X_0556_ u_buf.data\[2\]\[28\] _0141_ _0142_ i_instruction[28] _0152_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[28\] sky130_fd_sc_hs__a221o_1
X_0487_ _0111_ VSS VSS VCC VCC _0112_ sky130_fd_sc_hs__buf_2
X_1039_ clknet_4_5_0_i_clk u_buf.g_data\[2\].d_next\[12\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[12\] sky130_fd_sc_hs__dfxtp_1
X_1108_ clknet_4_6_0_i_clk u_buf.g_data\[0\].d_next\[15\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[15\] sky130_fd_sc_hs__dfxtp_1
X_0410_ o_pc[1] VSS VSS VCC VCC _0067_ sky130_fd_sc_hs__buf_2
X_0608_ u_buf.data\[1\]\[16\] _0178_ _0175_ i_instruction[16] _0184_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[16\] sky130_fd_sc_hs__a221o_1
X_0539_ u_buf.data\[3\]\[20\] _0143_ _0137_ VSS VSS VCC VCC _0144_ sky130_fd_sc_hs__and3_1
X_0890_ u_buf.data\[3\]\[27\] _0375_ _0376_ i_instruction[27] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[27\] sky130_fd_sc_hs__a22o_1
X_0873_ u_buf.data\[3\]\[12\] _0373_ _0374_ i_instruction[12] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[12\] sky130_fd_sc_hs__a22o_1
X_0942_ o_addr[11] _0338_ _0395_ VSS VSS VCC VCC _0035_ sky130_fd_sc_hs__mux2_1
X_1141_ clknet_4_2_0_i_clk _0017_ VSS VSS VCC VCC u_buf.latch_hi\[1\] sky130_fd_sc_hs__dfxtp_1
X_1072_ clknet_4_5_0_i_clk u_buf.g_data\[1\].d_next\[12\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[12\] sky130_fd_sc_hs__dfxtp_1
X_0787_ o_pc[7] _0302_ VSS VSS VCC VCC _0310_ sky130_fd_sc_hs__and2_1
X_0925_ o_addr[4] _0286_ _0395_ VSS VSS VCC VCC _0396_ sky130_fd_sc_hs__mux2_1
X_0856_ _0369_ VSS VSS VCC VCC _0370_ sky130_fd_sc_hs__buf_2
X_0641_ u_buf.data\[2\]\[31\] _0115_ _0157_ VSS VSS VCC VCC _0203_ sky130_fd_sc_hs__and3_1
X_0710_ u_buf.data\[1\]\[26\] _0235_ _0244_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[26\]
+ sky130_fd_sc_hs__a21o_1
X_0572_ _0158_ VSS VSS VCC VCC _0164_ sky130_fd_sc_hs__buf_2
X_1055_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[28\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[28\] sky130_fd_sc_hs__dfxtp_1
X_1124_ clknet_4_9_0_i_clk u_buf.g_data\[0\].d_next\[31\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[31\] sky130_fd_sc_hs__dfxtp_1
X_0839_ o_pc[13] _0343_ VSS VSS VCC VCC _0356_ sky130_fd_sc_hs__nand2_1
X_0908_ u_buf.is_head\[0\] u_buf.first_half VSS VSS VCC VCC o_ready sky130_fd_sc_hs__nor2_4
X_0624_ u_buf.data\[1\]\[22\] _0192_ _0189_ i_instruction[22] _0194_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[22\] sky130_fd_sc_hs__a221o_1
X_0555_ u_buf.data\[3\]\[28\] _0143_ _0114_ VSS VSS VCC VCC _0152_ sky130_fd_sc_hs__and3_1
X_0486_ _0110_ _0108_ VSS VSS VCC VCC _0111_ sky130_fd_sc_hs__nor2_1
X_1107_ clknet_4_6_0_i_clk u_buf.g_data\[0\].d_next\[14\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[14\] sky130_fd_sc_hs__dfxtp_1
X_1038_ clknet_4_5_0_i_clk u_buf.g_data\[2\].d_next\[11\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[11\] sky130_fd_sc_hs__dfxtp_1
X_0538_ _0110_ VSS VSS VCC VCC _0143_ sky130_fd_sc_hs__clkbuf_2
X_0607_ u_buf.data\[2\]\[16\] _0173_ _0176_ VSS VSS VCC VCC _0184_ sky130_fd_sc_hs__and3_1
X_0469_ _0098_ VSS VSS VCC VCC o_instruction[11] sky130_fd_sc_hs__buf_2
X_0941_ _0034_ VSS VSS VCC VCC _0010_ sky130_fd_sc_hs__clkbuf_1
X_0872_ u_buf.data\[3\]\[11\] _0373_ _0374_ i_instruction[11] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[11\] sky130_fd_sc_hs__a22o_1
X_1140_ clknet_4_0_0_i_clk _0016_ VSS VSS VCC VCC u_buf.latch_hi\[0\] sky130_fd_sc_hs__dfxtp_1
X_1071_ clknet_4_5_0_i_clk u_buf.g_data\[1\].d_next\[11\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[11\] sky130_fd_sc_hs__dfxtp_1
X_0924_ _0391_ VSS VSS VCC VCC _0395_ sky130_fd_sc_hs__inv_2
X_0786_ _0255_ i_pc_trap[7] _0308_ _0065_ VSS VSS VCC VCC _0309_ sky130_fd_sc_hs__o211a_1
X_0855_ _0114_ _0368_ VSS VSS VCC VCC _0369_ sky130_fd_sc_hs__nor2_2
X_0571_ i_instruction[0] _0160_ _0163_ VSS VSS VCC VCC u_buf.g_data\[1\].d_next\[0\]
+ sky130_fd_sc_hs__a21o_1
X_0640_ u_buf.data\[1\]\[30\] _0192_ _0159_ i_instruction[30] _0202_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[30\] sky130_fd_sc_hs__a221o_1
X_1123_ clknet_4_12_0_i_clk u_buf.g_data\[0\].d_next\[30\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[30\] sky130_fd_sc_hs__dfxtp_1
X_1054_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[27\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[27\] sky130_fd_sc_hs__dfxtp_1
X_0907_ _0386_ VSS VSS VCC VCC u_buf.g_data\[0\].h_next sky130_fd_sc_hs__clkbuf_1
X_0838_ o_pc[13] _0343_ VSS VSS VCC VCC _0355_ sky130_fd_sc_hs__or2_1
X_0769_ _0254_ i_pc_trap[5] _0292_ _0293_ i_reset_n VSS VSS VCC VCC _0294_
+ sky130_fd_sc_hs__o221a_1
X_0623_ u_buf.data\[2\]\[22\] _0187_ _0190_ VSS VSS VCC VCC _0194_ sky130_fd_sc_hs__and3_1
X_0554_ u_buf.data\[2\]\[27\] _0141_ _0142_ i_instruction[27] _0151_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[27\] sky130_fd_sc_hs__a221o_1
X_0485_ u_buf.is_head\[3\] _0105_ VSS VSS VCC VCC _0110_ sky130_fd_sc_hs__nor2_2
X_1106_ clknet_4_7_0_i_clk u_buf.g_data\[0\].d_next\[13\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[13\] sky130_fd_sc_hs__dfxtp_1
X_1037_ clknet_4_5_0_i_clk u_buf.g_data\[2\].d_next\[10\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[10\] sky130_fd_sc_hs__dfxtp_1
Xclkbuf_4_14_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_14_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0537_ _0111_ VSS VSS VCC VCC _0142_ sky130_fd_sc_hs__buf_2
X_0606_ u_buf.data\[1\]\[15\] _0178_ _0175_ i_instruction[15] _0183_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[15\] sky130_fd_sc_hs__a221o_1
X_0468_ u_buf.data\[0\]\[11\] u_buf.latch_hi\[11\] _0088_ VSS VSS VCC VCC
+ _0098_ sky130_fd_sc_hs__mux2_1
X_0940_ o_addr[10] _0331_ _0395_ VSS VSS VCC VCC _0034_ sky130_fd_sc_hs__mux2_1
X_0871_ u_buf.data\[3\]\[10\] _0373_ _0374_ i_instruction[10] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[10\] sky130_fd_sc_hs__a22o_1
X_1070_ clknet_4_4_0_i_clk u_buf.g_data\[1\].d_next\[10\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[10\] sky130_fd_sc_hs__dfxtp_1
X_0923_ _0394_ VSS VSS VCC VCC _0003_ sky130_fd_sc_hs__clkbuf_1
X_0854_ u_buf.is_head\[3\] u_buf.i_push _0104_ VSS VSS VCC VCC _0368_ sky130_fd_sc_hs__and3_1
X_0785_ _0256_ i_pc_target[7] _0305_ _0307_ i_ebreak VSS VSS VCC VCC _0308_
+ sky130_fd_sc_hs__a221o_1
X_0570_ u_buf.data\[2\]\[0\] _0161_ _0162_ _0158_ u_buf.data\[1\]\[0\] VSS VSS
+ VCC VCC _0163_ sky130_fd_sc_hs__a32o_1
X_1122_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[29\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[29\] sky130_fd_sc_hs__dfxtp_1
X_1053_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[26\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[26\] sky130_fd_sc_hs__dfxtp_1
X_0906_ _0251_ _0385_ VSS VSS VCC VCC _0386_ sky130_fd_sc_hs__and2_1
X_0837_ _0254_ i_pc_trap[13] _0352_ _0353_ i_reset_n VSS VSS VCC VCC _0354_
+ sky130_fd_sc_hs__o221a_1
X_0768_ _0270_ i_pc_target[5] _0258_ VSS VSS VCC VCC _0293_ sky130_fd_sc_hs__a21o_1
X_0699_ i_instruction[21] _0236_ _0237_ u_buf.data\[0\]\[21\] VSS VSS VCC VCC
+ _0239_ sky130_fd_sc_hs__a22o_1
Xclkbuf_4_10_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_10_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0553_ u_buf.data\[3\]\[27\] _0143_ _0114_ VSS VSS VCC VCC _0151_ sky130_fd_sc_hs__and3_1
X_0484_ _0108_ VSS VSS VCC VCC _0109_ sky130_fd_sc_hs__buf_2
X_0622_ u_buf.data\[1\]\[21\] _0192_ _0189_ i_instruction[21] _0193_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[21\] sky130_fd_sc_hs__a221o_1
X_1105_ clknet_4_4_0_i_clk u_buf.g_data\[0\].d_next\[12\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[12\] sky130_fd_sc_hs__dfxtp_1
X_1036_ clknet_4_6_0_i_clk u_buf.g_data\[2\].d_next\[9\] VSS VSS VCC VCC u_buf.data\[2\]\[9\]
+ sky130_fd_sc_hs__dfxtp_1
X_0605_ u_buf.data\[2\]\[15\] _0173_ _0176_ VSS VSS VCC VCC _0183_ sky130_fd_sc_hs__and3_1
X_0536_ _0108_ VSS VSS VCC VCC _0141_ sky130_fd_sc_hs__buf_2
X_0467_ _0097_ VSS VSS VCC VCC o_instruction[10] sky130_fd_sc_hs__buf_2
X_1019_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[25\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[25\] sky130_fd_sc_hs__dfxtp_1
X_0519_ u_buf.data\[3\]\[12\] _0129_ _0123_ VSS VSS VCC VCC _0132_ sky130_fd_sc_hs__and3_1
X_0870_ _0371_ VSS VSS VCC VCC _0374_ sky130_fd_sc_hs__buf_2
X_0999_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[5\] VSS VSS VCC VCC u_buf.data\[3\]\[5\]
+ sky130_fd_sc_hs__dfxtp_1
X_0853_ o_pc[15] _0252_ _0365_ _0264_ _0367_ VSS VSS VCC VCC o_pc_next[15]
+ sky130_fd_sc_hs__a221o_4
X_0922_ _0278_ o_addr[3] _0391_ VSS VSS VCC VCC _0394_ sky130_fd_sc_hs__mux2_1
X_0784_ _0256_ _0306_ VSS VSS VCC VCC _0307_ sky130_fd_sc_hs__nor2_1
X_1052_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[25\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[25\] sky130_fd_sc_hs__dfxtp_1
X_1121_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[28\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[28\] sky130_fd_sc_hs__dfxtp_1
X_0767_ _0257_ _0290_ _0291_ VSS VSS VCC VCC _0292_ sky130_fd_sc_hs__nor3_1
X_0905_ u_buf.is_head\[2\] _0378_ _0380_ u_buf.is_head\[1\] _0205_ VSS VSS VCC
+ VCC _0385_ sky130_fd_sc_hs__a221o_1
X_0836_ _0270_ i_pc_target[13] _0258_ VSS VSS VCC VCC _0353_ sky130_fd_sc_hs__a21o_1
X_0698_ u_buf.data\[1\]\[20\] _0235_ _0238_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[20\]
+ sky130_fd_sc_hs__a21o_1
X_0621_ u_buf.data\[2\]\[21\] _0187_ _0190_ VSS VSS VCC VCC _0193_ sky130_fd_sc_hs__and3_1
X_0552_ u_buf.data\[2\]\[26\] _0141_ _0142_ i_instruction[26] _0150_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[26\] sky130_fd_sc_hs__a221o_1
X_0483_ _0105_ _0107_ VSS VSS VCC VCC _0108_ sky130_fd_sc_hs__nor2_2
X_1035_ clknet_4_3_0_i_clk u_buf.g_data\[2\].d_next\[8\] VSS VSS VCC VCC u_buf.data\[2\]\[8\]
+ sky130_fd_sc_hs__dfxtp_1
X_1104_ clknet_4_4_0_i_clk u_buf.g_data\[0\].d_next\[11\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[11\] sky130_fd_sc_hs__dfxtp_1
X_0819_ _0254_ i_pc_trap[11] _0336_ _0337_ i_reset_n VSS VSS VCC VCC _0338_
+ sky130_fd_sc_hs__o221a_1
X_0604_ u_buf.data\[1\]\[14\] _0178_ _0175_ i_instruction[14] _0182_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[14\] sky130_fd_sc_hs__a221o_1
X_0535_ u_buf.data\[2\]\[19\] _0127_ _0128_ i_instruction[19] _0140_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[19\] sky130_fd_sc_hs__a221o_1
X_0466_ u_buf.data\[0\]\[10\] u_buf.latch_hi\[10\] _0088_ VSS VSS VCC VCC
+ _0097_ sky130_fd_sc_hs__mux2_1
Xclkbuf_4_8_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_8_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_1018_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[24\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[24\] sky130_fd_sc_hs__dfxtp_1
X_0518_ u_buf.data\[2\]\[11\] _0127_ _0128_ i_instruction[11] _0131_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[11\] sky130_fd_sc_hs__a221o_1
X_0449_ _0067_ VSS VSS VCC VCC _0088_ sky130_fd_sc_hs__clkbuf_4
X_0998_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[4\] VSS VSS VCC VCC u_buf.data\[3\]\[4\]
+ sky130_fd_sc_hs__dfxtp_1
X_0921_ _0393_ VSS VSS VCC VCC _0002_ sky130_fd_sc_hs__clkbuf_1
X_0852_ _0255_ i_pc_trap[15] _0366_ _0065_ VSS VSS VCC VCC _0367_ sky130_fd_sc_hs__o211a_1
X_0783_ o_addr[6] o_addr[7] _0290_ VSS VSS VCC VCC _0306_ sky130_fd_sc_hs__and3_1
X_1051_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[24\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[24\] sky130_fd_sc_hs__dfxtp_1
X_1120_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[27\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[27\] sky130_fd_sc_hs__dfxtp_1
X_0904_ _0377_ _0384_ VSS VSS VCC VCC u_buf.g_data\[1\].h_next sky130_fd_sc_hs__nor2_1
X_0766_ o_addr[5] _0283_ VSS VSS VCC VCC _0291_ sky130_fd_sc_hs__nor2_1
X_0835_ _0257_ _0350_ _0351_ VSS VSS VCC VCC _0352_ sky130_fd_sc_hs__nor3_1
X_0697_ i_instruction[20] _0236_ _0237_ u_buf.data\[0\]\[20\] VSS VSS VCC VCC
+ _0238_ sky130_fd_sc_hs__a22o_1
X_0551_ u_buf.data\[3\]\[26\] _0143_ _0137_ VSS VSS VCC VCC _0150_ sky130_fd_sc_hs__and3_1
X_0620_ _0158_ VSS VSS VCC VCC _0192_ sky130_fd_sc_hs__buf_2
X_0482_ u_buf.hi_valid _0106_ _0103_ VSS VSS VCC VCC _0107_ sky130_fd_sc_hs__a21oi_4
X_1034_ clknet_4_1_0_i_clk u_buf.g_data\[2\].d_next\[7\] VSS VSS VCC VCC u_buf.data\[2\]\[7\]
+ sky130_fd_sc_hs__dfxtp_1
X_1103_ clknet_4_5_0_i_clk u_buf.g_data\[0\].d_next\[10\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[10\] sky130_fd_sc_hs__dfxtp_1
Xclkbuf_4_4_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_4_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0749_ o_addr[2] o_addr[3] _0256_ VSS VSS VCC VCC _0276_ sky130_fd_sc_hs__o21ba_1
X_0818_ _0270_ i_pc_target[11] _0258_ VSS VSS VCC VCC _0337_ sky130_fd_sc_hs__a21o_1
X_0534_ u_buf.data\[3\]\[19\] _0129_ _0137_ VSS VSS VCC VCC _0140_ sky130_fd_sc_hs__and3_1
X_0603_ u_buf.data\[2\]\[14\] _0173_ _0176_ VSS VSS VCC VCC _0182_ sky130_fd_sc_hs__and3_1
X_0465_ _0096_ VSS VSS VCC VCC o_instruction[9] sky130_fd_sc_hs__buf_2
X_1017_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[23\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[23\] sky130_fd_sc_hs__dfxtp_1
X_0517_ u_buf.data\[3\]\[11\] _0129_ _0123_ VSS VSS VCC VCC _0131_ sky130_fd_sc_hs__and3_1
X_0448_ _0087_ VSS VSS VCC VCC o_instruction[1] sky130_fd_sc_hs__buf_2
X_0997_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[3\] VSS VSS VCC VCC u_buf.data\[3\]\[3\]
+ sky130_fd_sc_hs__dfxtp_1
X_0920_ _0273_ _0392_ _0391_ VSS VSS VCC VCC _0393_ sky130_fd_sc_hs__mux2_1
X_0782_ o_addr[6] _0290_ o_addr[7] VSS VSS VCC VCC _0305_ sky130_fd_sc_hs__a21o_1
X_0851_ _0257_ i_pc_target[15] _0258_ VSS VSS VCC VCC _0366_ sky130_fd_sc_hs__a21o_1
X_1050_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[23\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[23\] sky130_fd_sc_hs__dfxtp_1
X_0834_ o_addr[13] _0319_ _0349_ VSS VSS VCC VCC _0351_ sky130_fd_sc_hs__and3_1
X_0903_ u_buf.is_head\[2\] _0380_ _0383_ VSS VSS VCC VCC _0384_ sky130_fd_sc_hs__a21oi_1
X_0765_ o_addr[2] o_addr[3] o_addr[4] o_addr[5] VSS VSS VCC VCC _0290_ sky130_fd_sc_hs__and4_2
X_0696_ _0210_ VSS VSS VCC VCC _0237_ sky130_fd_sc_hs__buf_2
Xclkbuf_4_0_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_0_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0550_ u_buf.data\[2\]\[25\] _0141_ _0142_ i_instruction[25] _0149_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[25\] sky130_fd_sc_hs__a221o_1
X_0481_ u_buf.latch_hi\[0\] u_buf.latch_hi\[1\] _0067_ VSS VSS VCC VCC _0106_
+ sky130_fd_sc_hs__a21boi_4
X_1102_ clknet_4_3_0_i_clk u_buf.g_data\[0\].d_next\[9\] VSS VSS VCC VCC u_buf.data\[0\]\[9\]
+ sky130_fd_sc_hs__dfxtp_1
X_1033_ clknet_4_1_0_i_clk u_buf.g_data\[2\].d_next\[6\] VSS VSS VCC VCC u_buf.data\[2\]\[6\]
+ sky130_fd_sc_hs__dfxtp_1
X_0817_ _0257_ _0334_ _0335_ VSS VSS VCC VCC _0336_ sky130_fd_sc_hs__nor3_1
X_0748_ o_addr[2] o_addr[3] VSS VSS VCC VCC _0275_ sky130_fd_sc_hs__nand2_1
X_0679_ u_buf.data\[1\]\[12\] _0222_ _0227_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[12\]
+ sky130_fd_sc_hs__a21o_1
X_0533_ u_buf.data\[2\]\[18\] _0127_ _0128_ i_instruction[18] _0139_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[18\] sky130_fd_sc_hs__a221o_1
X_0602_ u_buf.data\[1\]\[13\] _0178_ _0175_ i_instruction[13] _0181_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[13\] sky130_fd_sc_hs__a221o_1
X_0464_ u_buf.data\[0\]\[9\] u_buf.latch_hi\[9\] _0088_ VSS VSS VCC VCC _0096_
+ sky130_fd_sc_hs__mux2_1
X_1016_ clknet_4_13_0_i_clk u_buf.g_data\[3\].d_next\[22\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[22\] sky130_fd_sc_hs__dfxtp_1
X_0516_ u_buf.data\[2\]\[10\] _0127_ _0128_ i_instruction[10] _0130_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[10\] sky130_fd_sc_hs__a221o_1
X_0447_ u_buf.data\[0\]\[1\] u_buf.latch_hi\[1\] _0077_ VSS VSS VCC VCC _0087_
+ sky130_fd_sc_hs__mux2_1
X_0996_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[2\] VSS VSS VCC VCC u_buf.data\[3\]\[2\]
+ sky130_fd_sc_hs__dfxtp_1
X_0850_ o_pc[15] _0362_ VSS VSS VCC VCC _0365_ sky130_fd_sc_hs__xor2_1
X_0781_ o_pc[6] _0253_ _0301_ o_pc_change _0304_ VSS VSS VCC VCC o_pc_next[6]
+ sky130_fd_sc_hs__a221o_4
X_0979_ _0056_ VSS VSS VCC VCC _0026_ sky130_fd_sc_hs__clkbuf_1
X_0902_ u_buf.is_head\[3\] _0378_ _0379_ u_buf.is_head\[1\] VSS VSS VCC VCC
+ _0383_ sky130_fd_sc_hs__a22o_1
X_0833_ _0319_ _0349_ o_addr[13] VSS VSS VCC VCC _0350_ sky130_fd_sc_hs__a21oi_1
X_0764_ o_pc[4] _0253_ _0286_ o_pc_change _0289_ VSS VSS VCC VCC o_pc_next[4]
+ sky130_fd_sc_hs__a221o_4
X_0695_ _0206_ VSS VSS VCC VCC _0236_ sky130_fd_sc_hs__buf_2
X_0480_ u_buf.i_push u_buf.is_head\[2\] _0104_ VSS VSS VCC VCC _0105_ sky130_fd_sc_hs__and3_1
X_1101_ clknet_4_2_0_i_clk u_buf.g_data\[0\].d_next\[8\] VSS VSS VCC VCC u_buf.data\[0\]\[8\]
+ sky130_fd_sc_hs__dfxtp_1
X_1032_ clknet_4_1_0_i_clk u_buf.g_data\[2\].d_next\[5\] VSS VSS VCC VCC u_buf.data\[2\]\[5\]
+ sky130_fd_sc_hs__dfxtp_1
X_0747_ o_pc[2] _0251_ _0268_ _0274_ VSS VSS VCC VCC o_pc_next[2] sky130_fd_sc_hs__a31o_4
X_0816_ o_addr[10] o_addr[11] _0319_ VSS VSS VCC VCC _0335_ sky130_fd_sc_hs__and3_1
X_0678_ i_instruction[12] _0223_ _0224_ u_buf.data\[0\]\[12\] VSS VSS VCC VCC
+ _0227_ sky130_fd_sc_hs__a22o_1
X_0601_ u_buf.data\[2\]\[13\] _0173_ _0176_ VSS VSS VCC VCC _0181_ sky130_fd_sc_hs__and3_1
X_0532_ u_buf.data\[3\]\[18\] _0129_ _0137_ VSS VSS VCC VCC _0139_ sky130_fd_sc_hs__and3_1
X_0463_ _0095_ VSS VSS VCC VCC o_instruction[8] sky130_fd_sc_hs__buf_2
X_1015_ clknet_4_13_0_i_clk u_buf.g_data\[3\].d_next\[21\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[21\] sky130_fd_sc_hs__dfxtp_1
X_0515_ u_buf.data\[3\]\[10\] _0129_ _0123_ VSS VSS VCC VCC _0130_ sky130_fd_sc_hs__and3_1
X_0446_ _0086_ VSS VSS VCC VCC o_instruction[0] sky130_fd_sc_hs__buf_2
X_0995_ clknet_4_6_0_i_clk u_buf.g_data\[3\].d_next\[1\] VSS VSS VCC VCC u_buf.data\[3\]\[1\]
+ sky130_fd_sc_hs__dfxtp_1
X_0429_ u_buf.data\[0\]\[24\] u_buf.data\[0\]\[8\] _0077_ VSS VSS VCC VCC
+ _0078_ sky130_fd_sc_hs__mux2_1
X_0780_ _0302_ _0303_ VSS VSS VCC VCC _0304_ sky130_fd_sc_hs__nor2_1
X_0978_ u_buf.data\[0\]\[26\] u_buf.latch_hi\[10\] _0250_ VSS VSS VCC VCC
+ _0056_ sky130_fd_sc_hs__mux2_1
X_0763_ _0287_ _0288_ _0263_ VSS VSS VCC VCC _0289_ sky130_fd_sc_hs__and3b_1
X_0832_ o_addr[10] o_addr[11] o_addr[12] VSS VSS VCC VCC _0349_ sky130_fd_sc_hs__and3_1
X_0901_ _0377_ _0382_ VSS VSS VCC VCC u_buf.g_data\[2\].h_next sky130_fd_sc_hs__nor2_1
X_0694_ _0207_ VSS VSS VCC VCC _0235_ sky130_fd_sc_hs__buf_2
X_1100_ clknet_4_2_0_i_clk u_buf.g_data\[0\].d_next\[7\] VSS VSS VCC VCC u_buf.data\[0\]\[7\]
+ sky130_fd_sc_hs__dfxtp_1
X_1031_ clknet_4_4_0_i_clk u_buf.g_data\[2\].d_next\[4\] VSS VSS VCC VCC u_buf.data\[2\]\[4\]
+ sky130_fd_sc_hs__dfxtp_1
X_0746_ _0269_ _0264_ _0267_ _0273_ _0064_ VSS VSS VCC VCC _0274_ sky130_fd_sc_hs__a32o_1
X_0815_ o_addr[10] _0319_ o_addr[11] VSS VSS VCC VCC _0334_ sky130_fd_sc_hs__a21oi_1
X_0677_ u_buf.data\[1\]\[11\] _0222_ _0226_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[11\]
+ sky130_fd_sc_hs__a21o_1
X_0531_ u_buf.data\[2\]\[17\] _0127_ _0128_ i_instruction[17] _0138_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[17\] sky130_fd_sc_hs__a221o_1
X_0600_ u_buf.data\[1\]\[12\] _0178_ _0175_ i_instruction[12] _0180_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[12\] sky130_fd_sc_hs__a221o_1
X_0462_ u_buf.data\[0\]\[8\] u_buf.latch_hi\[8\] _0088_ VSS VSS VCC VCC _0095_
+ sky130_fd_sc_hs__mux2_1
X_1014_ clknet_4_13_0_i_clk u_buf.g_data\[3\].d_next\[20\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[20\] sky130_fd_sc_hs__dfxtp_1
X_0729_ i_ebreak VSS VSS VCC VCC _0258_ sky130_fd_sc_hs__buf_2
X_0514_ _0110_ VSS VSS VCC VCC _0129_ sky130_fd_sc_hs__clkbuf_2
X_0445_ u_buf.data\[0\]\[0\] u_buf.latch_hi\[0\] _0077_ VSS VSS VCC VCC _0086_
+ sky130_fd_sc_hs__mux2_1
X_0994_ clknet_4_6_0_i_clk u_buf.g_data\[3\].d_next\[0\] VSS VSS VCC VCC u_buf.data\[3\]\[0\]
+ sky130_fd_sc_hs__dfxtp_1
X_0428_ _0067_ VSS VSS VCC VCC _0077_ sky130_fd_sc_hs__clkbuf_4
X_0977_ _0055_ VSS VSS VCC VCC _0025_ sky130_fd_sc_hs__clkbuf_1
X_0900_ u_buf.is_head\[3\] _0380_ _0381_ VSS VSS VCC VCC _0382_ sky130_fd_sc_hs__a21oi_1
X_0831_ o_pc[12] _0253_ _0345_ _0348_ VSS VSS VCC VCC o_pc_next[12] sky130_fd_sc_hs__a211o_4
X_0762_ o_pc[2] o_pc[3] _0267_ o_pc[4] VSS VSS VCC VCC _0288_ sky130_fd_sc_hs__a31o_1
X_0693_ u_buf.data\[1\]\[19\] _0222_ _0234_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[19\]
+ sky130_fd_sc_hs__a21o_1
X_1030_ clknet_4_1_0_i_clk u_buf.g_data\[2\].d_next\[3\] VSS VSS VCC VCC u_buf.data\[2\]\[3\]
+ sky130_fd_sc_hs__dfxtp_1
X_0814_ o_pc[10] _0253_ _0331_ o_pc_change _0333_ VSS VSS VCC VCC o_pc_next[10]
+ sky130_fd_sc_hs__a221o_4
X_0745_ _0254_ i_pc_trap[2] _0272_ i_reset_n VSS VSS VCC VCC _0273_ sky130_fd_sc_hs__o211a_1
X_0676_ i_instruction[11] _0223_ _0224_ u_buf.data\[0\]\[11\] VSS VSS VCC VCC
+ _0226_ sky130_fd_sc_hs__a22o_1
X_1159_ clknet_4_8_0_i_clk o_pc_next[3] VSS VSS VCC VCC o_pc[3] sky130_fd_sc_hs__dfxtp_4
X_0530_ u_buf.data\[3\]\[17\] _0129_ _0137_ VSS VSS VCC VCC _0138_ sky130_fd_sc_hs__and3_1
X_0461_ _0094_ VSS VSS VCC VCC o_instruction[7] sky130_fd_sc_hs__buf_2
X_1013_ clknet_4_13_0_i_clk u_buf.g_data\[3\].d_next\[19\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[19\] sky130_fd_sc_hs__dfxtp_1
X_0728_ _0256_ VSS VSS VCC VCC _0257_ sky130_fd_sc_hs__buf_2
X_0659_ i_instruction[4] _0209_ _0211_ u_buf.data\[0\]\[4\] VSS VSS VCC VCC
+ _0216_ sky130_fd_sc_hs__a22o_1
X_0513_ _0111_ VSS VSS VCC VCC _0128_ sky130_fd_sc_hs__buf_2
X_0444_ _0085_ VSS VSS VCC VCC o_instruction[31] sky130_fd_sc_hs__buf_2
X_0993_ clknet_4_9_0_i_clk u_buf.g_data\[3\].h_next VSS VSS VCC VCC u_buf.is_head\[4\]
+ sky130_fd_sc_hs__dfxtp_1
X_0427_ _0076_ VSS VSS VCC VCC o_instruction[23] sky130_fd_sc_hs__buf_2
X_0976_ u_buf.data\[0\]\[25\] u_buf.latch_hi\[9\] _0045_ VSS VSS VCC VCC _0055_
+ sky130_fd_sc_hs__mux2_1
X_0830_ _0346_ _0347_ VSS VSS VCC VCC _0348_ sky130_fd_sc_hs__nor2_1
X_0761_ o_pc[2] o_pc[3] o_pc[4] _0267_ VSS VSS VCC VCC _0287_ sky130_fd_sc_hs__and4_1
X_0692_ i_instruction[19] _0223_ _0224_ u_buf.data\[0\]\[19\] VSS VSS VCC VCC
+ _0234_ sky130_fd_sc_hs__a22o_1
X_0959_ _0046_ VSS VSS VCC VCC _0016_ sky130_fd_sc_hs__clkbuf_1
X_0813_ o_pc[10] _0325_ _0332_ VSS VSS VCC VCC _0333_ sky130_fd_sc_hs__o21a_1
X_0744_ _0270_ i_pc_target[2] _0271_ _0258_ VSS VSS VCC VCC _0272_ sky130_fd_sc_hs__a211o_1
X_0675_ u_buf.data\[1\]\[10\] _0222_ _0225_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[10\]
+ sky130_fd_sc_hs__a21o_1
X_1158_ clknet_4_8_0_i_clk o_pc_next[2] VSS VSS VCC VCC o_pc[2] sky130_fd_sc_hs__dfxtp_4
X_1089_ clknet_4_14_0_i_clk u_buf.g_data\[1\].d_next\[29\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[29\] sky130_fd_sc_hs__dfxtp_1
X_0460_ u_buf.data\[0\]\[7\] u_buf.latch_hi\[7\] _0088_ VSS VSS VCC VCC _0094_
+ sky130_fd_sc_hs__mux2_1
X_1012_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[18\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[18\] sky130_fd_sc_hs__dfxtp_1
X_0727_ i_pc_select VSS VSS VCC VCC _0256_ sky130_fd_sc_hs__buf_2
X_0658_ u_buf.data\[1\]\[3\] _0208_ _0215_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[3\]
+ sky130_fd_sc_hs__a21o_1
X_0589_ _0114_ VSS VSS VCC VCC _0173_ sky130_fd_sc_hs__clkbuf_2
X_0512_ _0108_ VSS VSS VCC VCC _0127_ sky130_fd_sc_hs__buf_2
X_0443_ u_buf.data\[0\]\[31\] u_buf.data\[0\]\[15\] _0077_ VSS VSS VCC VCC
+ _0085_ sky130_fd_sc_hs__mux2_1
X_0992_ clknet_4_9_0_i_clk u_buf.is_head_next_0 VSS VSS VCC VCC u_buf.is_head\[0\]
+ sky130_fd_sc_hs__dfxtp_1
X_0426_ u_buf.data\[0\]\[23\] u_buf.data\[0\]\[7\] _0068_ VSS VSS VCC VCC
+ _0076_ sky130_fd_sc_hs__mux2_1
X_0975_ _0054_ VSS VSS VCC VCC _0024_ sky130_fd_sc_hs__clkbuf_1
X_0409_ _0066_ VSS VSS VCC VCC push_next sky130_fd_sc_hs__clkbuf_1
X_0760_ _0255_ i_pc_trap[4] _0285_ _0065_ VSS VSS VCC VCC _0286_ sky130_fd_sc_hs__o211a_1
X_0691_ u_buf.data\[1\]\[18\] _0222_ _0233_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[18\]
+ sky130_fd_sc_hs__a21o_1
X_0889_ u_buf.data\[3\]\[26\] _0375_ _0376_ i_instruction[26] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[26\] sky130_fd_sc_hs__a22o_1
X_0958_ u_buf.data\[0\]\[16\] u_buf.latch_hi\[0\] _0045_ VSS VSS VCC VCC _0046_
+ sky130_fd_sc_hs__mux2_1
X_0812_ o_pc[10] _0325_ _0263_ VSS VSS VCC VCC _0332_ sky130_fd_sc_hs__a21boi_1
X_0743_ _0256_ o_addr[2] VSS VSS VCC VCC _0271_ sky130_fd_sc_hs__nor2_1
X_0674_ i_instruction[10] _0223_ _0224_ u_buf.data\[0\]\[10\] VSS VSS VCC VCC
+ _0225_ sky130_fd_sc_hs__a22o_1
X_1157_ clknet_4_8_0_i_clk o_pc_next[1] VSS VSS VCC VCC o_pc[1] sky130_fd_sc_hs__dfxtp_2
X_1088_ clknet_4_14_0_i_clk u_buf.g_data\[1\].d_next\[28\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[28\] sky130_fd_sc_hs__dfxtp_1
X_1011_ clknet_4_7_0_i_clk u_buf.g_data\[3\].d_next\[17\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[17\] sky130_fd_sc_hs__dfxtp_1
X_0726_ _0254_ VSS VSS VCC VCC _0255_ sky130_fd_sc_hs__buf_2
X_0657_ i_instruction[3] _0209_ _0211_ u_buf.data\[0\]\[3\] VSS VSS VCC VCC
+ _0215_ sky130_fd_sc_hs__a22o_1
X_0588_ u_buf.data\[1\]\[8\] _0164_ _0160_ i_instruction[8] _0172_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[8\] sky130_fd_sc_hs__a221o_1
X_0511_ u_buf.data\[2\]\[9\] _0109_ _0112_ i_instruction[9] _0126_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[9\] sky130_fd_sc_hs__a221o_1
Xclkbuf_4_13_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_13_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0442_ _0084_ VSS VSS VCC VCC o_instruction[30] sky130_fd_sc_hs__buf_2
X_0709_ i_instruction[26] _0236_ _0237_ u_buf.data\[0\]\[26\] VSS VSS VCC VCC
+ _0244_ sky130_fd_sc_hs__a22o_1
X_0991_ _0377_ _0062_ VSS VSS VCC VCC _0032_ sky130_fd_sc_hs__nor2_1
X_0425_ _0075_ VSS VSS VCC VCC o_instruction[22] sky130_fd_sc_hs__buf_2
X_0974_ u_buf.data\[0\]\[24\] u_buf.latch_hi\[8\] _0045_ VSS VSS VCC VCC _0054_
+ sky130_fd_sc_hs__mux2_1
X_0408_ _0065_ i_ack _0063_ VSS VSS VCC VCC _0066_ sky130_fd_sc_hs__and3_1
X_0690_ i_instruction[18] _0223_ _0224_ u_buf.data\[0\]\[18\] VSS VSS VCC VCC
+ _0233_ sky130_fd_sc_hs__a22o_1
X_1173_ clknet_4_9_0_i_clk push_next VSS VSS VCC VCC u_buf.i_push sky130_fd_sc_hs__dfxtp_2
X_0888_ u_buf.data\[3\]\[25\] _0375_ _0376_ i_instruction[25] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[25\] sky130_fd_sc_hs__a22o_1
X_0957_ _0250_ VSS VSS VCC VCC _0045_ sky130_fd_sc_hs__clkbuf_4
X_0811_ _0254_ i_pc_trap[10] _0330_ i_reset_n VSS VSS VCC VCC _0331_ sky130_fd_sc_hs__o211a_1
X_0742_ _0256_ VSS VSS VCC VCC _0270_ sky130_fd_sc_hs__buf_2
X_0673_ _0210_ VSS VSS VCC VCC _0224_ sky130_fd_sc_hs__buf_2
X_1156_ clknet_4_8_0_i_clk _0000_ VSS VSS VCC VCC u_buf.first_half sky130_fd_sc_hs__dfxtp_1
X_1087_ clknet_4_14_0_i_clk u_buf.g_data\[1\].d_next\[27\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[27\] sky130_fd_sc_hs__dfxtp_1
X_1010_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[16\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[16\] sky130_fd_sc_hs__dfxtp_1
X_0725_ i_ebreak VSS VSS VCC VCC _0254_ sky130_fd_sc_hs__clkinv_2
X_0656_ u_buf.data\[1\]\[2\] _0208_ _0214_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[2\]
+ sky130_fd_sc_hs__a21o_1
X_0587_ u_buf.data\[2\]\[8\] _0161_ _0162_ VSS VSS VCC VCC _0172_ sky130_fd_sc_hs__and3_1
X_1139_ clknet_4_11_0_i_clk _0015_ VSS VSS VCC VCC o_addr[15] sky130_fd_sc_hs__dfxtp_4
X_0510_ u_buf.data\[3\]\[9\] _0113_ _0123_ VSS VSS VCC VCC _0126_ sky130_fd_sc_hs__and3_1
X_0441_ u_buf.data\[0\]\[30\] u_buf.data\[0\]\[14\] _0077_ VSS VSS VCC VCC
+ _0084_ sky130_fd_sc_hs__mux2_1
X_0639_ u_buf.data\[2\]\[30\] _0115_ _0157_ VSS VSS VCC VCC _0202_ sky130_fd_sc_hs__and3_1
X_0708_ u_buf.data\[1\]\[25\] _0235_ _0243_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[25\]
+ sky130_fd_sc_hs__a21o_1
X_0990_ u_buf.i_push _0262_ u_buf.hi_valid VSS VSS VCC VCC _0062_ sky130_fd_sc_hs__a21oi_1
X_0424_ u_buf.data\[0\]\[22\] u_buf.data\[0\]\[6\] _0068_ VSS VSS VCC VCC
+ _0075_ sky130_fd_sc_hs__mux2_1
X_0973_ _0053_ VSS VSS VCC VCC _0023_ sky130_fd_sc_hs__clkbuf_1
X_0407_ i_reset_n VSS VSS VCC VCC _0065_ sky130_fd_sc_hs__buf_2
X_1172_ clknet_4_8_0_i_clk _0032_ VSS VSS VCC VCC u_buf.hi_valid sky130_fd_sc_hs__dfxtp_1
X_0956_ o_addr[15] _0391_ _0043_ _0044_ VSS VSS VCC VCC _0015_ sky130_fd_sc_hs__a22o_1
X_0887_ u_buf.data\[3\]\[24\] _0375_ _0376_ i_instruction[24] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[24\] sky130_fd_sc_hs__a22o_1
X_0810_ _0256_ i_pc_target[10] _0328_ _0329_ i_ebreak VSS VSS VCC VCC _0330_
+ sky130_fd_sc_hs__a221o_1
X_0741_ o_pc[2] VSS VSS VCC VCC _0269_ sky130_fd_sc_hs__inv_2
X_0672_ _0206_ VSS VSS VCC VCC _0223_ sky130_fd_sc_hs__buf_2
X_1155_ clknet_4_8_0_i_clk _0031_ VSS VSS VCC VCC u_buf.latch_hi\[15\] sky130_fd_sc_hs__dfxtp_1
X_1086_ clknet_4_15_0_i_clk u_buf.g_data\[1\].d_next\[26\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[26\] sky130_fd_sc_hs__dfxtp_1
X_0939_ _0033_ VSS VSS VCC VCC _0009_ sky130_fd_sc_hs__clkbuf_1
X_0724_ _0252_ VSS VSS VCC VCC _0253_ sky130_fd_sc_hs__buf_4
X_0655_ i_instruction[2] _0209_ _0211_ u_buf.data\[0\]\[2\] VSS VSS VCC VCC
+ _0214_ sky130_fd_sc_hs__a22o_1
X_0586_ u_buf.data\[1\]\[7\] _0164_ _0160_ i_instruction[7] _0171_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[7\] sky130_fd_sc_hs__a221o_1
X_1069_ clknet_4_3_0_i_clk u_buf.g_data\[1\].d_next\[9\] VSS VSS VCC VCC u_buf.data\[1\]\[9\]
+ sky130_fd_sc_hs__dfxtp_1
X_1138_ clknet_4_11_0_i_clk _0014_ VSS VSS VCC VCC o_addr[14] sky130_fd_sc_hs__dfxtp_4
X_0440_ _0083_ VSS VSS VCC VCC o_instruction[29] sky130_fd_sc_hs__buf_2
X_0707_ i_instruction[25] _0236_ _0237_ u_buf.data\[0\]\[25\] VSS VSS VCC VCC
+ _0243_ sky130_fd_sc_hs__a22o_1
Xclkbuf_4_7_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_7_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0569_ _0157_ VSS VSS VCC VCC _0162_ sky130_fd_sc_hs__clkbuf_2
X_0638_ u_buf.data\[1\]\[29\] _0192_ _0189_ i_instruction[29] _0201_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[29\] sky130_fd_sc_hs__a221o_1
X_0423_ _0074_ VSS VSS VCC VCC o_instruction[21] sky130_fd_sc_hs__buf_2
X_0972_ u_buf.data\[0\]\[23\] u_buf.latch_hi\[7\] _0045_ VSS VSS VCC VCC _0053_
+ sky130_fd_sc_hs__mux2_1
X_0406_ _0064_ VSS VSS VCC VCC o_pc_change sky130_fd_sc_hs__buf_4
X_1171_ clknet_4_10_0_i_clk o_pc_next[15] VSS VSS VCC VCC o_pc[15] sky130_fd_sc_hs__dfxtp_4
X_0886_ u_buf.data\[3\]\[23\] _0375_ _0376_ i_instruction[23] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[23\] sky130_fd_sc_hs__a22o_1
X_0955_ _0255_ i_pc_trap[15] _0395_ _0065_ VSS VSS VCC VCC _0044_ sky130_fd_sc_hs__o211a_1
X_0740_ u_buf.first_half _0250_ _0267_ VSS VSS VCC VCC _0268_ sky130_fd_sc_hs__or3b_1
X_0671_ _0207_ VSS VSS VCC VCC _0222_ sky130_fd_sc_hs__buf_2
X_1154_ clknet_4_2_0_i_clk _0030_ VSS VSS VCC VCC u_buf.latch_hi\[14\] sky130_fd_sc_hs__dfxtp_1
X_1085_ clknet_4_14_0_i_clk u_buf.g_data\[1\].d_next\[25\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[25\] sky130_fd_sc_hs__dfxtp_1
X_0869_ _0369_ VSS VSS VCC VCC _0373_ sky130_fd_sc_hs__buf_2
X_0938_ o_addr[9] _0323_ _0395_ VSS VSS VCC VCC _0033_ sky130_fd_sc_hs__mux2_1
X_0723_ u_buf.first_half _0250_ _0251_ VSS VSS VCC VCC _0252_ sky130_fd_sc_hs__o21a_2
X_0654_ u_buf.data\[1\]\[1\] _0208_ _0213_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[1\]
+ sky130_fd_sc_hs__a21o_1
X_0585_ u_buf.data\[2\]\[7\] _0161_ _0162_ VSS VSS VCC VCC _0171_ sky130_fd_sc_hs__and3_1
Xclkbuf_4_3_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_3_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_1137_ clknet_4_11_0_i_clk _0013_ VSS VSS VCC VCC o_addr[13] sky130_fd_sc_hs__dfxtp_4
X_1068_ clknet_4_3_0_i_clk u_buf.g_data\[1\].d_next\[8\] VSS VSS VCC VCC u_buf.data\[1\]\[8\]
+ sky130_fd_sc_hs__dfxtp_1
X_0706_ u_buf.data\[1\]\[24\] _0235_ _0242_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[24\]
+ sky130_fd_sc_hs__a21o_1
X_0568_ _0107_ VSS VSS VCC VCC _0161_ sky130_fd_sc_hs__clkbuf_2
X_0499_ u_buf.data\[3\]\[4\] _0113_ _0115_ VSS VSS VCC VCC _0120_ sky130_fd_sc_hs__and3_1
X_0637_ u_buf.data\[2\]\[29\] _0115_ _0190_ VSS VSS VCC VCC _0201_ sky130_fd_sc_hs__and3_1
X_0422_ u_buf.data\[0\]\[21\] u_buf.data\[0\]\[5\] _0068_ VSS VSS VCC VCC
+ _0074_ sky130_fd_sc_hs__mux2_1
X_0971_ _0052_ VSS VSS VCC VCC _0022_ sky130_fd_sc_hs__clkbuf_1
X_0405_ _0063_ VSS VSS VCC VCC _0064_ sky130_fd_sc_hs__inv_2
X_1170_ clknet_4_10_0_i_clk o_pc_next[14] VSS VSS VCC VCC o_pc[14] sky130_fd_sc_hs__dfxtp_4
X_0885_ u_buf.data\[3\]\[22\] _0375_ _0376_ i_instruction[22] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[22\] sky130_fd_sc_hs__a22o_1
X_0954_ _0041_ _0042_ _0366_ VSS VSS VCC VCC _0043_ sky130_fd_sc_hs__a21o_1
X_0670_ u_buf.data\[1\]\[9\] _0208_ _0221_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[9\]
+ sky130_fd_sc_hs__a21o_1
X_1153_ clknet_4_2_0_i_clk _0029_ VSS VSS VCC VCC u_buf.latch_hi\[13\] sky130_fd_sc_hs__dfxtp_1
X_1084_ clknet_4_14_0_i_clk u_buf.g_data\[1\].d_next\[24\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[24\] sky130_fd_sc_hs__dfxtp_1
X_0799_ o_addr[6] _0290_ _0317_ o_addr[9] VSS VSS VCC VCC _0320_ sky130_fd_sc_hs__a31o_1
X_0937_ o_addr[8] _0391_ _0402_ _0403_ VSS VSS VCC VCC _0008_ sky130_fd_sc_hs__a22o_1
X_0868_ u_buf.data\[3\]\[9\] _0370_ _0372_ i_instruction[9] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[9\] sky130_fd_sc_hs__a22o_1
X_0722_ i_reset_n _0063_ VSS VSS VCC VCC _0251_ sky130_fd_sc_hs__and2_1
X_0653_ i_instruction[1] _0209_ _0211_ u_buf.data\[0\]\[1\] VSS VSS VCC VCC
+ _0213_ sky130_fd_sc_hs__a22o_1
X_0584_ u_buf.data\[1\]\[6\] _0164_ _0160_ i_instruction[6] _0170_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[6\] sky130_fd_sc_hs__a221o_1
X_1136_ clknet_4_11_0_i_clk _0012_ VSS VSS VCC VCC o_addr[12] sky130_fd_sc_hs__dfxtp_2
X_1067_ clknet_4_1_0_i_clk u_buf.g_data\[1\].d_next\[7\] VSS VSS VCC VCC u_buf.data\[1\]\[7\]
+ sky130_fd_sc_hs__dfxtp_1
X_0705_ i_instruction[24] _0236_ _0237_ u_buf.data\[0\]\[24\] VSS VSS VCC VCC
+ _0242_ sky130_fd_sc_hs__a22o_1
X_0636_ u_buf.data\[1\]\[28\] _0192_ _0189_ i_instruction[28] _0200_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[28\] sky130_fd_sc_hs__a221o_1
X_0567_ _0159_ VSS VSS VCC VCC _0160_ sky130_fd_sc_hs__buf_2
X_0498_ u_buf.data\[2\]\[3\] _0109_ _0112_ i_instruction[3] _0119_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[3\] sky130_fd_sc_hs__a221o_1
X_1119_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[26\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[26\] sky130_fd_sc_hs__dfxtp_1
X_0421_ _0073_ VSS VSS VCC VCC o_instruction[20] sky130_fd_sc_hs__buf_2
X_0619_ u_buf.data\[1\]\[20\] _0178_ _0189_ i_instruction[20] _0191_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[20\] sky130_fd_sc_hs__a221o_1
X_0970_ u_buf.data\[0\]\[22\] u_buf.latch_hi\[6\] _0045_ VSS VSS VCC VCC _0052_
+ sky130_fd_sc_hs__mux2_1
X_0404_ i_ebreak i_pc_select VSS VSS VCC VCC _0063_ sky130_fd_sc_hs__nor2_1
X_0884_ u_buf.data\[3\]\[21\] _0375_ _0376_ i_instruction[21] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[21\] sky130_fd_sc_hs__a22o_1
X_0953_ o_addr[14] o_addr[15] _0351_ _0257_ VSS VSS VCC VCC _0042_ sky130_fd_sc_hs__a31oi_1
X_1152_ clknet_4_2_0_i_clk _0028_ VSS VSS VCC VCC u_buf.latch_hi\[12\] sky130_fd_sc_hs__dfxtp_1
X_1083_ clknet_4_15_0_i_clk u_buf.g_data\[1\].d_next\[23\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[23\] sky130_fd_sc_hs__dfxtp_1
X_0936_ _0314_ _0391_ VSS VSS VCC VCC _0403_ sky130_fd_sc_hs__nor2_1
X_0798_ _0318_ VSS VSS VCC VCC _0319_ sky130_fd_sc_hs__clkbuf_2
X_0867_ u_buf.data\[3\]\[8\] _0370_ _0372_ i_instruction[8] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[8\] sky130_fd_sc_hs__a22o_1
X_0721_ _0103_ VSS VSS VCC VCC _0250_ sky130_fd_sc_hs__clkbuf_4
X_0652_ u_buf.data\[1\]\[0\] _0208_ _0212_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[0\]
+ sky130_fd_sc_hs__a21o_1
X_0583_ u_buf.data\[2\]\[6\] _0161_ _0162_ VSS VSS VCC VCC _0170_ sky130_fd_sc_hs__and3_1
X_1135_ clknet_4_10_0_i_clk _0011_ VSS VSS VCC VCC o_addr[11] sky130_fd_sc_hs__dfxtp_4
X_1066_ clknet_4_3_0_i_clk u_buf.g_data\[1\].d_next\[6\] VSS VSS VCC VCC u_buf.data\[1\]\[6\]
+ sky130_fd_sc_hs__dfxtp_1
X_0919_ _0255_ i_pc_trap[2] _0272_ VSS VSS VCC VCC _0392_ sky130_fd_sc_hs__o21ai_1
X_0566_ _0157_ _0158_ VSS VSS VCC VCC _0159_ sky130_fd_sc_hs__nor2_1
X_0704_ u_buf.data\[1\]\[23\] _0235_ _0241_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[23\]
+ sky130_fd_sc_hs__a21o_1
X_0635_ u_buf.data\[2\]\[28\] _0187_ _0190_ VSS VSS VCC VCC _0200_ sky130_fd_sc_hs__and3_1
X_0497_ u_buf.data\[3\]\[3\] _0113_ _0115_ VSS VSS VCC VCC _0119_ sky130_fd_sc_hs__and3_1
X_1049_ clknet_4_13_0_i_clk u_buf.g_data\[2\].d_next\[22\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[22\] sky130_fd_sc_hs__dfxtp_1
X_1118_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[25\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[25\] sky130_fd_sc_hs__dfxtp_1
X_0420_ u_buf.data\[0\]\[20\] u_buf.data\[0\]\[4\] _0068_ VSS VSS VCC VCC
+ _0073_ sky130_fd_sc_hs__mux2_1
X_0549_ u_buf.data\[3\]\[25\] _0143_ _0137_ VSS VSS VCC VCC _0149_ sky130_fd_sc_hs__and3_1
X_0618_ u_buf.data\[2\]\[20\] _0187_ _0190_ VSS VSS VCC VCC _0191_ sky130_fd_sc_hs__and3_1
X_0952_ o_addr[14] _0351_ o_addr[15] VSS VSS VCC VCC _0041_ sky130_fd_sc_hs__a21o_1
X_0883_ u_buf.data\[3\]\[20\] _0375_ _0376_ i_instruction[20] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[20\] sky130_fd_sc_hs__a22o_1
X_1151_ clknet_4_2_0_i_clk _0027_ VSS VSS VCC VCC u_buf.latch_hi\[11\] sky130_fd_sc_hs__dfxtp_1
X_1082_ clknet_4_13_0_i_clk u_buf.g_data\[1\].d_next\[22\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[22\] sky130_fd_sc_hs__dfxtp_1
X_0935_ _0257_ _0401_ _0315_ VSS VSS VCC VCC _0402_ sky130_fd_sc_hs__o21ai_1
X_0866_ u_buf.data\[3\]\[7\] _0370_ _0372_ i_instruction[7] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[7\] sky130_fd_sc_hs__a22o_1
X_0797_ o_addr[6] o_addr[9] _0290_ _0317_ VSS VSS VCC VCC _0318_ sky130_fd_sc_hs__and4_1
X_0720_ u_buf.data\[1\]\[31\] _0207_ _0249_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[31\]
+ sky130_fd_sc_hs__a21o_1
X_0582_ u_buf.data\[1\]\[5\] _0164_ _0160_ i_instruction[5] _0169_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[5\] sky130_fd_sc_hs__a221o_1
X_0651_ i_instruction[0] _0209_ _0211_ u_buf.data\[0\]\[0\] VSS VSS VCC VCC
+ _0212_ sky130_fd_sc_hs__a22o_1
X_1134_ clknet_4_11_0_i_clk _0010_ VSS VSS VCC VCC o_addr[10] sky130_fd_sc_hs__dfxtp_4
X_1065_ clknet_4_1_0_i_clk u_buf.g_data\[1\].d_next\[5\] VSS VSS VCC VCC u_buf.data\[1\]\[5\]
+ sky130_fd_sc_hs__dfxtp_1
X_0849_ o_pc[14] _0252_ _0361_ _0064_ _0364_ VSS VSS VCC VCC o_pc_next[14]
+ sky130_fd_sc_hs__a221o_4
X_0918_ o_addr[1] _0391_ _0260_ VSS VSS VCC VCC _0001_ sky130_fd_sc_hs__a21o_1
X_0703_ i_instruction[23] _0236_ _0237_ u_buf.data\[0\]\[23\] VSS VSS VCC VCC
+ _0241_ sky130_fd_sc_hs__a22o_1
X_0565_ _0107_ _0156_ VSS VSS VCC VCC _0158_ sky130_fd_sc_hs__nor2_2
X_0496_ u_buf.data\[2\]\[2\] _0109_ _0112_ i_instruction[2] _0118_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[2\] sky130_fd_sc_hs__a221o_1
X_0634_ u_buf.data\[1\]\[27\] _0192_ _0189_ i_instruction[27] _0199_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[27\] sky130_fd_sc_hs__a221o_1
X_1117_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[24\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[24\] sky130_fd_sc_hs__dfxtp_1
X_1048_ clknet_4_13_0_i_clk u_buf.g_data\[2\].d_next\[21\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[21\] sky130_fd_sc_hs__dfxtp_1
X_0548_ u_buf.data\[2\]\[24\] _0141_ _0142_ i_instruction[24] _0148_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[24\] sky130_fd_sc_hs__a221o_1
X_0479_ _0067_ _0103_ VSS VSS VCC VCC _0104_ sky130_fd_sc_hs__or2_1
X_0617_ _0157_ VSS VSS VCC VCC _0190_ sky130_fd_sc_hs__clkbuf_2
X_0882_ _0371_ VSS VSS VCC VCC _0376_ sky130_fd_sc_hs__buf_2
X_0951_ _0040_ VSS VSS VCC VCC _0014_ sky130_fd_sc_hs__clkbuf_1
X_1150_ clknet_4_2_0_i_clk _0026_ VSS VSS VCC VCC u_buf.latch_hi\[10\] sky130_fd_sc_hs__dfxtp_1
X_1081_ clknet_4_13_0_i_clk u_buf.g_data\[1\].d_next\[21\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[21\] sky130_fd_sc_hs__dfxtp_1
X_0934_ o_addr[6] _0290_ _0317_ _0400_ VSS VSS VCC VCC _0401_ sky130_fd_sc_hs__a31o_1
X_0865_ u_buf.data\[3\]\[6\] _0370_ _0372_ i_instruction[6] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[6\] sky130_fd_sc_hs__a22o_1
X_0796_ o_addr[7] o_addr[8] VSS VSS VCC VCC _0317_ sky130_fd_sc_hs__and2_1
X_0650_ _0210_ VSS VSS VCC VCC _0211_ sky130_fd_sc_hs__buf_2
X_0581_ u_buf.data\[2\]\[5\] _0161_ _0162_ VSS VSS VCC VCC _0169_ sky130_fd_sc_hs__and3_1
X_1064_ clknet_4_1_0_i_clk u_buf.g_data\[1\].d_next\[4\] VSS VSS VCC VCC u_buf.data\[1\]\[4\]
+ sky130_fd_sc_hs__dfxtp_1
X_1133_ clknet_4_11_0_i_clk _0009_ VSS VSS VCC VCC o_addr[9] sky130_fd_sc_hs__dfxtp_2
X_0848_ _0362_ _0263_ _0363_ VSS VSS VCC VCC _0364_ sky130_fd_sc_hs__and3b_1
X_0779_ o_pc[6] _0295_ _0264_ VSS VSS VCC VCC _0303_ sky130_fd_sc_hs__o21ai_1
X_0917_ i_ack o_cyc _0377_ VSS VSS VCC VCC _0391_ sky130_fd_sc_hs__a21oi_4
X_0702_ u_buf.data\[1\]\[22\] _0235_ _0240_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[22\]
+ sky130_fd_sc_hs__a21o_1
X_0633_ u_buf.data\[2\]\[27\] _0187_ _0190_ VSS VSS VCC VCC _0199_ sky130_fd_sc_hs__and3_1
X_0564_ u_buf.is_head\[2\] _0156_ VSS VSS VCC VCC _0157_ sky130_fd_sc_hs__nor2_2
X_0495_ u_buf.data\[3\]\[2\] _0113_ _0115_ VSS VSS VCC VCC _0118_ sky130_fd_sc_hs__and3_1
X_1047_ clknet_4_13_0_i_clk u_buf.g_data\[2\].d_next\[20\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[20\] sky130_fd_sc_hs__dfxtp_1
X_1116_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[23\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[23\] sky130_fd_sc_hs__dfxtp_1
X_0616_ _0159_ VSS VSS VCC VCC _0189_ sky130_fd_sc_hs__buf_2
X_0547_ u_buf.data\[3\]\[24\] _0143_ _0137_ VSS VSS VCC VCC _0148_ sky130_fd_sc_hs__and3_1
X_0478_ u_buf.is_head\[0\] i_stall VSS VSS VCC VCC _0103_ sky130_fd_sc_hs__or2_2
X_0881_ _0369_ VSS VSS VCC VCC _0375_ sky130_fd_sc_hs__buf_2
X_0950_ o_addr[14] _0361_ _0395_ VSS VSS VCC VCC _0040_ sky130_fd_sc_hs__mux2_1
X_1080_ clknet_4_13_0_i_clk u_buf.g_data\[1\].d_next\[20\] VSS VSS VCC VCC
+ u_buf.data\[1\]\[20\] sky130_fd_sc_hs__dfxtp_1
X_0795_ o_pc[8] _0253_ _0313_ _0264_ _0316_ VSS VSS VCC VCC o_pc_next[8] sky130_fd_sc_hs__a221o_4
X_0933_ o_addr[8] _0306_ VSS VSS VCC VCC _0400_ sky130_fd_sc_hs__nor2_1
X_0864_ u_buf.data\[3\]\[5\] _0370_ _0372_ i_instruction[5] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[5\] sky130_fd_sc_hs__a22o_1
X_0580_ u_buf.data\[1\]\[4\] _0164_ _0160_ i_instruction[4] _0168_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[4\] sky130_fd_sc_hs__a221o_1
X_1063_ clknet_4_1_0_i_clk u_buf.g_data\[1\].d_next\[3\] VSS VSS VCC VCC u_buf.data\[1\]\[3\]
+ sky130_fd_sc_hs__dfxtp_1
X_1132_ clknet_4_11_0_i_clk _0008_ VSS VSS VCC VCC o_addr[8] sky130_fd_sc_hs__dfxtp_4
X_0916_ _0390_ VSS VSS VCC VCC u_buf.g_data\[3\].h_next sky130_fd_sc_hs__clkbuf_1
X_0847_ o_pc[13] _0343_ o_pc[14] VSS VSS VCC VCC _0363_ sky130_fd_sc_hs__a21o_1
X_0778_ o_pc[5] o_pc[6] _0287_ VSS VSS VCC VCC _0302_ sky130_fd_sc_hs__and3_1
X_0563_ u_buf.i_push u_buf.is_head\[1\] _0104_ VSS VSS VCC VCC _0156_ sky130_fd_sc_hs__and3_1
X_0701_ i_instruction[22] _0236_ _0237_ u_buf.data\[0\]\[22\] VSS VSS VCC VCC
+ _0240_ sky130_fd_sc_hs__a22o_1
X_0632_ u_buf.data\[1\]\[26\] _0192_ _0189_ i_instruction[26] _0198_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[26\] sky130_fd_sc_hs__a221o_1
X_0494_ u_buf.data\[2\]\[1\] _0109_ _0112_ i_instruction[1] _0117_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[1\] sky130_fd_sc_hs__a221o_1
X_1046_ clknet_4_13_0_i_clk u_buf.g_data\[2\].d_next\[19\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[19\] sky130_fd_sc_hs__dfxtp_1
X_1115_ clknet_4_12_0_i_clk u_buf.g_data\[0\].d_next\[22\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[22\] sky130_fd_sc_hs__dfxtp_1
X_0546_ u_buf.data\[2\]\[23\] _0141_ _0142_ i_instruction[23] _0147_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[23\] sky130_fd_sc_hs__a221o_1
X_0615_ u_buf.data\[1\]\[19\] _0178_ _0175_ i_instruction[19] _0188_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[19\] sky130_fd_sc_hs__a221o_1
X_0477_ _0102_ VSS VSS VCC VCC o_instruction[15] sky130_fd_sc_hs__buf_2
X_1029_ clknet_4_1_0_i_clk u_buf.g_data\[2\].d_next\[2\] VSS VSS VCC VCC u_buf.data\[2\]\[2\]
+ sky130_fd_sc_hs__dfxtp_1
X_0529_ _0107_ VSS VSS VCC VCC _0137_ sky130_fd_sc_hs__clkbuf_2
X_0880_ u_buf.data\[3\]\[19\] _0373_ _0374_ i_instruction[19] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[19\] sky130_fd_sc_hs__a22o_1
X_0932_ _0399_ VSS VSS VCC VCC _0007_ sky130_fd_sc_hs__clkbuf_1
X_0794_ _0314_ _0315_ VSS VSS VCC VCC _0316_ sky130_fd_sc_hs__nor2_1
X_0863_ u_buf.data\[3\]\[4\] _0370_ _0372_ i_instruction[4] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[4\] sky130_fd_sc_hs__a22o_1
X_1131_ clknet_4_11_0_i_clk _0007_ VSS VSS VCC VCC o_addr[7] sky130_fd_sc_hs__dfxtp_4
X_1062_ clknet_4_1_0_i_clk u_buf.g_data\[1\].d_next\[2\] VSS VSS VCC VCC u_buf.data\[1\]\[2\]
+ sky130_fd_sc_hs__dfxtp_1
X_0915_ _0251_ _0389_ VSS VSS VCC VCC _0390_ sky130_fd_sc_hs__and2_1
X_0846_ o_pc[13] o_pc[14] _0343_ VSS VSS VCC VCC _0362_ sky130_fd_sc_hs__and3_1
X_0777_ _0255_ i_pc_trap[6] _0300_ _0065_ VSS VSS VCC VCC _0301_ sky130_fd_sc_hs__o211a_1
X_0700_ u_buf.data\[1\]\[21\] _0235_ _0239_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[21\]
+ sky130_fd_sc_hs__a21o_1
X_0562_ u_buf.data\[2\]\[31\] _0108_ _0111_ i_instruction[31] _0155_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[31\] sky130_fd_sc_hs__a221o_1
X_0631_ u_buf.data\[2\]\[26\] _0187_ _0190_ VSS VSS VCC VCC _0198_ sky130_fd_sc_hs__and3_1
X_0493_ u_buf.data\[3\]\[1\] _0113_ _0115_ VSS VSS VCC VCC _0117_ sky130_fd_sc_hs__and3_1
X_1114_ clknet_4_12_0_i_clk u_buf.g_data\[0\].d_next\[21\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[21\] sky130_fd_sc_hs__dfxtp_1
X_1045_ clknet_4_7_0_i_clk u_buf.g_data\[2\].d_next\[18\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[18\] sky130_fd_sc_hs__dfxtp_1
X_0829_ _0257_ i_pc_target[12] _0258_ VSS VSS VCC VCC _0347_ sky130_fd_sc_hs__a21oi_1
Xclkbuf_4_12_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_12_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0545_ u_buf.data\[3\]\[23\] _0143_ _0137_ VSS VSS VCC VCC _0147_ sky130_fd_sc_hs__and3_1
X_0476_ u_buf.data\[0\]\[15\] u_buf.latch_hi\[15\] _0067_ VSS VSS VCC VCC
+ _0102_ sky130_fd_sc_hs__mux2_1
X_0614_ u_buf.data\[2\]\[19\] _0187_ _0176_ VSS VSS VCC VCC _0188_ sky130_fd_sc_hs__and3_1
X_1028_ clknet_4_3_0_i_clk u_buf.g_data\[2\].d_next\[1\] VSS VSS VCC VCC u_buf.data\[2\]\[1\]
+ sky130_fd_sc_hs__dfxtp_1
X_0528_ u_buf.data\[2\]\[16\] _0127_ _0128_ i_instruction[16] _0136_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[16\] sky130_fd_sc_hs__a221o_1
X_0459_ _0093_ VSS VSS VCC VCC o_instruction[6] sky130_fd_sc_hs__buf_2
X_0931_ o_addr[7] _0309_ _0395_ VSS VSS VCC VCC _0399_ sky130_fd_sc_hs__mux2_1
X_0862_ u_buf.data\[3\]\[3\] _0370_ _0372_ i_instruction[3] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[3\] sky130_fd_sc_hs__a22o_1
X_0793_ _0257_ i_pc_target[8] _0258_ VSS VSS VCC VCC _0315_ sky130_fd_sc_hs__a21oi_1
X_1130_ clknet_4_10_0_i_clk _0006_ VSS VSS VCC VCC o_addr[6] sky130_fd_sc_hs__dfxtp_4
X_1061_ clknet_4_3_0_i_clk u_buf.g_data\[1\].d_next\[1\] VSS VSS VCC VCC u_buf.data\[1\]\[1\]
+ sky130_fd_sc_hs__dfxtp_1
X_0914_ u_buf.is_head\[3\] _0379_ _0380_ u_buf.is_head\[4\] VSS VSS VCC VCC
+ _0389_ sky130_fd_sc_hs__a22o_1
X_0845_ _0254_ i_pc_trap[14] _0359_ _0360_ i_reset_n VSS VSS VCC VCC _0361_
+ sky130_fd_sc_hs__o221a_1
X_0776_ _0270_ i_pc_target[6] _0298_ _0299_ i_ebreak VSS VSS VCC VCC _0300_
+ sky130_fd_sc_hs__a221o_1
X_0492_ u_buf.data\[2\]\[0\] _0109_ _0112_ i_instruction[0] _0116_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[0\] sky130_fd_sc_hs__a221o_1
X_0561_ u_buf.data\[3\]\[31\] _0110_ _0114_ VSS VSS VCC VCC _0155_ sky130_fd_sc_hs__and3_1
X_0630_ u_buf.data\[1\]\[25\] _0192_ _0189_ i_instruction[25] _0197_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[25\] sky130_fd_sc_hs__a221o_1
X_1044_ clknet_4_7_0_i_clk u_buf.g_data\[2\].d_next\[17\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[17\] sky130_fd_sc_hs__dfxtp_1
X_1113_ clknet_4_12_0_i_clk u_buf.g_data\[0\].d_next\[20\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[20\] sky130_fd_sc_hs__dfxtp_1
X_0828_ _0255_ i_pc_trap[12] _0065_ VSS VSS VCC VCC _0346_ sky130_fd_sc_hs__o21ai_1
X_0759_ _0270_ i_pc_target[4] _0282_ _0284_ i_ebreak VSS VSS VCC VCC _0285_
+ sky130_fd_sc_hs__a221o_1
X_0613_ _0114_ VSS VSS VCC VCC _0187_ sky130_fd_sc_hs__clkbuf_2
X_0544_ u_buf.data\[2\]\[22\] _0141_ _0142_ i_instruction[22] _0146_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[22\] sky130_fd_sc_hs__a221o_1
X_0475_ _0101_ VSS VSS VCC VCC o_instruction[14] sky130_fd_sc_hs__buf_2
X_1027_ clknet_4_3_0_i_clk u_buf.g_data\[2\].d_next\[0\] VSS VSS VCC VCC u_buf.data\[2\]\[0\]
+ sky130_fd_sc_hs__dfxtp_1
X_0527_ u_buf.data\[3\]\[16\] _0129_ _0123_ VSS VSS VCC VCC _0136_ sky130_fd_sc_hs__and3_1
X_0458_ u_buf.data\[0\]\[6\] u_buf.latch_hi\[6\] _0088_ VSS VSS VCC VCC _0093_
+ sky130_fd_sc_hs__mux2_1
X_0930_ _0398_ VSS VSS VCC VCC _0006_ sky130_fd_sc_hs__clkbuf_1
X_0792_ _0255_ i_pc_trap[8] _0065_ VSS VSS VCC VCC _0314_ sky130_fd_sc_hs__o21ai_1
X_0861_ u_buf.data\[3\]\[2\] _0370_ _0372_ i_instruction[2] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[2\] sky130_fd_sc_hs__a22o_1
X_1060_ clknet_4_3_0_i_clk u_buf.g_data\[1\].d_next\[0\] VSS VSS VCC VCC u_buf.data\[1\]\[0\]
+ sky130_fd_sc_hs__dfxtp_1
X_0913_ u_buf.is_head\[3\] u_buf.i_push _0103_ u_buf.is_head\[4\] VSS VSS VCC
+ VCC o_cyc sky130_fd_sc_hs__a31oi_4
X_0775_ o_addr[6] _0290_ _0256_ VSS VSS VCC VCC _0299_ sky130_fd_sc_hs__o21ba_1
X_0844_ _0270_ i_pc_target[14] _0258_ VSS VSS VCC VCC _0360_ sky130_fd_sc_hs__a21o_1
X_0491_ u_buf.data\[3\]\[0\] _0113_ _0115_ VSS VSS VCC VCC _0116_ sky130_fd_sc_hs__and3_1
X_0560_ u_buf.data\[2\]\[30\] _0108_ _0111_ i_instruction[30] _0154_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[30\] sky130_fd_sc_hs__a221o_1
X_1043_ clknet_4_5_0_i_clk u_buf.g_data\[2\].d_next\[16\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[16\] sky130_fd_sc_hs__dfxtp_1
X_1112_ clknet_4_6_0_i_clk u_buf.g_data\[0\].d_next\[19\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[19\] sky130_fd_sc_hs__dfxtp_1
X_0827_ _0343_ _0344_ _0264_ VSS VSS VCC VCC _0345_ sky130_fd_sc_hs__and3b_1
X_0758_ _0256_ _0283_ VSS VSS VCC VCC _0284_ sky130_fd_sc_hs__nor2_1
X_0689_ u_buf.data\[1\]\[17\] _0222_ _0232_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[17\]
+ sky130_fd_sc_hs__a21o_1
X_0612_ u_buf.data\[1\]\[18\] _0178_ _0175_ i_instruction[18] _0186_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[18\] sky130_fd_sc_hs__a221o_1
X_0543_ u_buf.data\[3\]\[22\] _0143_ _0137_ VSS VSS VCC VCC _0146_ sky130_fd_sc_hs__and3_1
X_0474_ u_buf.data\[0\]\[14\] u_buf.latch_hi\[14\] _0067_ VSS VSS VCC VCC
+ _0101_ sky130_fd_sc_hs__mux2_1
X_1026_ clknet_4_9_0_i_clk u_buf.g_data\[2\].h_next VSS VSS VCC VCC u_buf.is_head\[3\]
+ sky130_fd_sc_hs__dfxtp_2
Xclkbuf_4_6_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_6_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0526_ u_buf.data\[2\]\[15\] _0127_ _0128_ i_instruction[15] _0135_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[15\] sky130_fd_sc_hs__a221o_1
X_0457_ _0092_ VSS VSS VCC VCC o_instruction[5] sky130_fd_sc_hs__buf_2
X_1009_ clknet_4_7_0_i_clk u_buf.g_data\[3\].d_next\[15\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[15\] sky130_fd_sc_hs__dfxtp_1
X_0509_ u_buf.data\[2\]\[8\] _0109_ _0112_ i_instruction[8] _0125_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[8\] sky130_fd_sc_hs__a221o_1
X_0791_ o_pc[8] _0310_ VSS VSS VCC VCC _0313_ sky130_fd_sc_hs__xor2_1
X_0860_ u_buf.data\[3\]\[1\] _0370_ _0372_ i_instruction[1] VSS VSS VCC VCC
+ u_buf.g_data\[3\].d_next\[1\] sky130_fd_sc_hs__a22o_1
X_0989_ _0061_ VSS VSS VCC VCC _0031_ sky130_fd_sc_hs__clkbuf_1
X_0912_ u_buf.i_push _0388_ _0251_ VSS VSS VCC VCC u_buf.is_head_next_0 sky130_fd_sc_hs__o21ai_1
X_0774_ o_addr[6] _0290_ VSS VSS VCC VCC _0298_ sky130_fd_sc_hs__nand2_1
X_0843_ o_addr[14] _0351_ _0358_ VSS VSS VCC VCC _0359_ sky130_fd_sc_hs__o21ba_1
X_0490_ _0114_ VSS VSS VCC VCC _0115_ sky130_fd_sc_hs__clkbuf_2
X_1042_ clknet_4_7_0_i_clk u_buf.g_data\[2\].d_next\[15\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[15\] sky130_fd_sc_hs__dfxtp_1
X_1111_ clknet_4_7_0_i_clk u_buf.g_data\[0\].d_next\[18\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[18\] sky130_fd_sc_hs__dfxtp_1
X_0826_ o_pc[10] o_pc[11] _0325_ o_pc[12] VSS VSS VCC VCC _0344_ sky130_fd_sc_hs__a31o_1
X_0757_ o_addr[2] o_addr[3] o_addr[4] VSS VSS VCC VCC _0283_ sky130_fd_sc_hs__and3_1
Xclkbuf_4_2_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_4_2_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0688_ i_instruction[17] _0223_ _0224_ u_buf.data\[0\]\[17\] VSS VSS VCC VCC
+ _0232_ sky130_fd_sc_hs__a22o_1
X_0611_ u_buf.data\[2\]\[18\] _0173_ _0176_ VSS VSS VCC VCC _0186_ sky130_fd_sc_hs__and3_1
X_0542_ u_buf.data\[2\]\[21\] _0141_ _0142_ i_instruction[21] _0145_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[21\] sky130_fd_sc_hs__a221o_1
X_0473_ _0100_ VSS VSS VCC VCC o_instruction[13] sky130_fd_sc_hs__buf_2
X_1025_ clknet_4_6_0_i_clk u_buf.g_data\[3\].d_next\[31\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[31\] sky130_fd_sc_hs__dfxtp_1
X_0809_ o_addr[10] _0319_ i_pc_select VSS VSS VCC VCC _0329_ sky130_fd_sc_hs__o21ba_1
X_0525_ u_buf.data\[3\]\[15\] _0129_ _0123_ VSS VSS VCC VCC _0135_ sky130_fd_sc_hs__and3_1
X_0456_ u_buf.data\[0\]\[5\] u_buf.latch_hi\[5\] _0088_ VSS VSS VCC VCC _0092_
+ sky130_fd_sc_hs__mux2_1
X_1008_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[14\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[14\] sky130_fd_sc_hs__dfxtp_1
X_0439_ u_buf.data\[0\]\[29\] u_buf.data\[0\]\[13\] _0077_ VSS VSS VCC VCC
+ _0083_ sky130_fd_sc_hs__mux2_1
X_0508_ u_buf.data\[3\]\[8\] _0113_ _0123_ VSS VSS VCC VCC _0125_ sky130_fd_sc_hs__and3_1
X_0790_ o_pc[7] _0253_ _0309_ o_pc_change _0312_ VSS VSS VCC VCC o_pc_next[7]
+ sky130_fd_sc_hs__a221o_4
X_0988_ u_buf.data\[0\]\[31\] u_buf.latch_hi\[15\] _0250_ VSS VSS VCC VCC
+ _0061_ sky130_fd_sc_hs__mux2_1
X_0911_ u_buf.is_head\[1\] _0161_ u_buf.is_head\[0\] VSS VSS VCC VCC _0388_
+ sky130_fd_sc_hs__a21oi_1
X_0842_ o_addr[13] o_addr[14] _0319_ _0349_ _0256_ VSS VSS VCC VCC _0358_
+ sky130_fd_sc_hs__a41o_1
X_0773_ o_pc[5] _0253_ _0294_ o_pc_change _0297_ VSS VSS VCC VCC o_pc_next[5]
+ sky130_fd_sc_hs__a221o_4
X_1110_ clknet_4_6_0_i_clk u_buf.g_data\[0\].d_next\[17\] VSS VSS VCC VCC
+ u_buf.data\[0\]\[17\] sky130_fd_sc_hs__dfxtp_1
X_1041_ clknet_4_5_0_i_clk u_buf.g_data\[2\].d_next\[14\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[14\] sky130_fd_sc_hs__dfxtp_1
X_0825_ o_pc[5] _0287_ _0324_ _0342_ VSS VSS VCC VCC _0343_ sky130_fd_sc_hs__and4_1
X_0756_ o_addr[2] o_addr[3] o_addr[4] VSS VSS VCC VCC _0282_ sky130_fd_sc_hs__a21o_1
X_0687_ u_buf.data\[1\]\[16\] _0222_ _0231_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[16\]
+ sky130_fd_sc_hs__a21o_1
X_0541_ u_buf.data\[3\]\[21\] _0143_ _0137_ VSS VSS VCC VCC _0145_ sky130_fd_sc_hs__and3_1
X_0610_ u_buf.data\[1\]\[17\] _0178_ _0175_ i_instruction[17] _0185_ VSS VSS VCC
+ VCC u_buf.g_data\[1\].d_next\[17\] sky130_fd_sc_hs__a221o_1
X_0472_ u_buf.data\[0\]\[13\] u_buf.latch_hi\[13\] _0067_ VSS VSS VCC VCC
+ _0100_ sky130_fd_sc_hs__mux2_1
X_1024_ clknet_4_12_0_i_clk u_buf.g_data\[3\].d_next\[30\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[30\] sky130_fd_sc_hs__dfxtp_1
X_0808_ o_addr[10] _0319_ VSS VSS VCC VCC _0328_ sky130_fd_sc_hs__nand2_1
X_0739_ u_buf.data\[0\]\[0\] u_buf.data\[0\]\[1\] o_pc[1] VSS VSS VCC VCC
+ _0267_ sky130_fd_sc_hs__a21o_1
X_0524_ u_buf.data\[2\]\[14\] _0127_ _0128_ i_instruction[14] _0134_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[14\] sky130_fd_sc_hs__a221o_1
X_0455_ _0091_ VSS VSS VCC VCC o_instruction[4] sky130_fd_sc_hs__buf_2
X_1007_ clknet_4_7_0_i_clk u_buf.g_data\[3\].d_next\[13\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[13\] sky130_fd_sc_hs__dfxtp_1
X_0438_ _0082_ VSS VSS VCC VCC o_instruction[28] sky130_fd_sc_hs__buf_2
X_0507_ u_buf.data\[2\]\[7\] _0109_ _0112_ i_instruction[7] _0124_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[7\] sky130_fd_sc_hs__a221o_1
X_0987_ _0060_ VSS VSS VCC VCC _0030_ sky130_fd_sc_hs__clkbuf_1
X_0841_ o_pc[13] _0252_ _0354_ o_pc_change _0357_ VSS VSS VCC VCC o_pc_next[13]
+ sky130_fd_sc_hs__a221o_4
X_0772_ _0295_ _0296_ VSS VSS VCC VCC _0297_ sky130_fd_sc_hs__nor2_1
X_0910_ _0387_ VSS VSS VCC VCC _0000_ sky130_fd_sc_hs__clkbuf_1
X_1040_ clknet_4_7_0_i_clk u_buf.g_data\[2\].d_next\[13\] VSS VSS VCC VCC
+ u_buf.data\[2\]\[13\] sky130_fd_sc_hs__dfxtp_1
X_0755_ o_pc[3] _0253_ _0278_ o_pc_change _0281_ VSS VSS VCC VCC o_pc_next[3]
+ sky130_fd_sc_hs__a221o_4
X_0824_ o_pc[9] o_pc[10] o_pc[11] o_pc[12] VSS VSS VCC VCC _0342_ sky130_fd_sc_hs__and4_1
X_0686_ i_instruction[16] _0223_ _0224_ u_buf.data\[0\]\[16\] VSS VSS VCC VCC
+ _0231_ sky130_fd_sc_hs__a22o_1
X_1169_ clknet_4_10_0_i_clk o_pc_next[13] VSS VSS VCC VCC o_pc[13] sky130_fd_sc_hs__dfxtp_4
X_0540_ u_buf.data\[2\]\[20\] _0141_ _0142_ i_instruction[20] _0144_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[20\] sky130_fd_sc_hs__a221o_1
X_0471_ _0099_ VSS VSS VCC VCC o_instruction[12] sky130_fd_sc_hs__buf_2
X_1023_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[29\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[29\] sky130_fd_sc_hs__dfxtp_1
X_0738_ _0068_ _0253_ _0260_ _0266_ VSS VSS VCC VCC o_pc_next[1] sky130_fd_sc_hs__a211o_4
X_0807_ o_pc[9] _0253_ _0323_ o_pc_change _0327_ VSS VSS VCC VCC o_pc_next[9]
+ sky130_fd_sc_hs__a221o_4
X_0669_ i_instruction[9] _0209_ _0211_ u_buf.data\[0\]\[9\] VSS VSS VCC VCC
+ _0221_ sky130_fd_sc_hs__a22o_1
X_0523_ u_buf.data\[3\]\[14\] _0129_ _0123_ VSS VSS VCC VCC _0134_ sky130_fd_sc_hs__and3_1
X_0454_ u_buf.data\[0\]\[4\] u_buf.latch_hi\[4\] _0088_ VSS VSS VCC VCC _0091_
+ sky130_fd_sc_hs__mux2_1
X_1006_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[12\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[12\] sky130_fd_sc_hs__dfxtp_1
X_0506_ u_buf.data\[3\]\[7\] _0113_ _0123_ VSS VSS VCC VCC _0124_ sky130_fd_sc_hs__and3_1
X_0437_ u_buf.data\[0\]\[28\] u_buf.data\[0\]\[12\] _0077_ VSS VSS VCC VCC
+ _0082_ sky130_fd_sc_hs__mux2_1
X_0986_ u_buf.data\[0\]\[30\] u_buf.latch_hi\[14\] _0250_ VSS VSS VCC VCC
+ _0060_ sky130_fd_sc_hs__mux2_1
X_0840_ _0263_ _0355_ _0356_ VSS VSS VCC VCC _0357_ sky130_fd_sc_hs__and3_1
X_0771_ o_pc[5] _0287_ _0264_ VSS VSS VCC VCC _0296_ sky130_fd_sc_hs__o21ai_1
X_0969_ _0051_ VSS VSS VCC VCC _0021_ sky130_fd_sc_hs__clkbuf_1
X_0754_ _0264_ _0279_ _0280_ VSS VSS VCC VCC _0281_ sky130_fd_sc_hs__and3_1
X_0823_ o_pc[11] _0252_ _0338_ o_pc_change _0341_ VSS VSS VCC VCC o_pc_next[11]
+ sky130_fd_sc_hs__a221o_4
X_0685_ u_buf.data\[1\]\[15\] _0222_ _0230_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[15\]
+ sky130_fd_sc_hs__a21o_1
X_1168_ clknet_4_10_0_i_clk o_pc_next[12] VSS VSS VCC VCC o_pc[12] sky130_fd_sc_hs__dfxtp_4
X_1099_ clknet_4_0_0_i_clk u_buf.g_data\[0\].d_next\[6\] VSS VSS VCC VCC u_buf.data\[0\]\[6\]
+ sky130_fd_sc_hs__dfxtp_1
X_0470_ u_buf.data\[0\]\[12\] u_buf.latch_hi\[12\] _0067_ VSS VSS VCC VCC
+ _0099_ sky130_fd_sc_hs__mux2_1
X_1022_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[28\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[28\] sky130_fd_sc_hs__dfxtp_1
X_0737_ _0067_ _0261_ _0264_ _0265_ VSS VSS VCC VCC _0266_ sky130_fd_sc_hs__o211a_1
X_0806_ _0325_ _0263_ _0326_ VSS VSS VCC VCC _0327_ sky130_fd_sc_hs__and3b_1
X_0668_ u_buf.data\[1\]\[8\] _0208_ _0220_ VSS VSS VCC VCC u_buf.g_data\[0\].d_next\[8\]
+ sky130_fd_sc_hs__a21o_1
X_0599_ u_buf.data\[2\]\[12\] _0173_ _0176_ VSS VSS VCC VCC _0180_ sky130_fd_sc_hs__and3_1
X_0522_ u_buf.data\[2\]\[13\] _0127_ _0128_ i_instruction[13] _0133_ VSS VSS VCC
+ VCC u_buf.g_data\[2\].d_next\[13\] sky130_fd_sc_hs__a221o_1
X_0453_ _0090_ VSS VSS VCC VCC o_instruction[3] sky130_fd_sc_hs__buf_2
X_1005_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[11\] VSS VSS VCC VCC
+ u_buf.data\[3\]\[11\] sky130_fd_sc_hs__dfxtp_1
X_0505_ _0107_ VSS VSS VCC VCC _0123_ sky130_fd_sc_hs__clkbuf_2
X_0436_ _0081_ VSS VSS VCC VCC o_instruction[27] sky130_fd_sc_hs__buf_2
