
.include ../../elements/inc_lib.spice
.include simulation/rom.spice

.param VCC=1.8

VVCC VCC 0 PWL 0ns 0 1ns 0 1.1ns {VCC}
VVSS VSS 0 PWL 0n 0

.include simulation/stimuli_rom.cir

.OPTIONS MEASURE MEASFAIL=1
*.OPTIONS LINSOL type=AztecOO AZ_tol=1.0e-3 TR_PARTITION=1
.OPTIONS TIMEINT RELTOL=1e-3 ABSTOL=1e-5 method=gear
.OPTIONS DIST STRATEGY=2

.tran 1p 200n
.print tran format=raw file=simulation/rom.spice.raw v(*) i(*)

*.meas tran rd_v_0[*] find v(rd[*]) at=1.8n

.meas tran power avg par('(-1*v(VCC)*I(VVCC))') from=1.4n to=19n

.GLOBAL VCC
.GLOBAL VSS
.end
