* NGSPICE file created from rv_ctrl.ext - technology: sky130A


X_66_ clknet_1_0__leaf_i_clk _00_ VSS VSS VCC VCC inst_sup\[0\] sky130_fd_sc_hd__dfxtp_2
X_49_ i_alu1_rd[1] i_alu1_rd[0] i_alu1_rd[3] i_alu1_rd[4] VSS VSS VCC VCC
+ _20_ sky130_fd_sc_hd__nor4_1
X_65_ inst_sup\[0\] _23_ o_alu2_flush _29_ VSS VSS VCC VCC _01_ sky130_fd_sc_hd__a211o_2
X_48_ _13_ _14_ _15_ _18_ VSS VSS VCC VCC _19_ sky130_fd_sc_hd__or4_1
X_64_ o_alu1_stall i_need_pause _22_ inst_sup\[1\] VSS VSS VCC VCC _29_ sky130_fd_sc_hd__o31a_1
X_47_ _04_ i_decode_rs2[1] _16_ i_alu1_rd[2] _17_ VSS VSS VCC VCC _18_ sky130_fd_sc_hd__a221o_1
X_63_ i_decode_inst_sup _23_ o_alu2_flush _28_ VSS VSS VCC VCC _00_ sky130_fd_sc_hd__a211o_2
X_46_ i_alu1_rd[4] i_decode_rs2[4] VSS VSS VCC VCC _17_ sky130_fd_sc_hd__xor2_1
X_62_ o_alu1_stall i_need_pause _22_ inst_sup\[0\] VSS VSS VCC VCC _28_ sky130_fd_sc_hd__o31a_1
X_45_ i_decode_rs2[2] VSS VSS VCC VCC _16_ sky130_fd_sc_hd__inv_2
Xclkbuf_0_i_clk i_clk VSS VSS VCC VCC clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_61_ _27_ VSS VSS VCC VCC o_write_flush sky130_fd_sc_hd__buf_2
X_44_ _04_ i_decode_rs2[1] i_decode_rs2[2] _02_ VSS VSS VCC VCC _15_ sky130_fd_sc_hd__a2bb2o_1
X_60_ o_alu1_stall o_alu2_flush VSS VSS VCC VCC _27_ sky130_fd_sc_hd__or2_1
X_43_ i_alu1_rd[3] i_decode_rs2[3] VSS VSS VCC VCC _14_ sky130_fd_sc_hd__xor2_1
X_42_ i_alu1_rd[0] i_decode_rs2[0] VSS VSS VCC VCC _13_ sky130_fd_sc_hd__xor2_1
X_41_ _03_ _05_ _09_ _11_ VSS VSS VCC VCC _12_ sky130_fd_sc_hd__or4b_1
X_40_ _06_ i_decode_rs1[3] i_decode_rs1[4] _07_ _10_ VSS VSS VCC VCC _11_
+ sky130_fd_sc_hd__o221a_1
X_59_ _26_ VSS VSS VCC VCC o_alu1_flush sky130_fd_sc_hd__buf_2
X_58_ o_alu2_flush _25_ VSS VSS VCC VCC _26_ sky130_fd_sc_hd__or2_1
X_57_ i_need_pause _22_ i_alu2_ready VSS VSS VCC VCC _25_ sky130_fd_sc_hd__o21a_1
X_56_ _24_ VSS VSS VCC VCC o_alu2_flush sky130_fd_sc_hd__clkbuf_4
X_39_ i_decode_rs1[1] i_alu1_rd[1] VSS VSS VCC VCC _10_ sky130_fd_sc_hd__or2b_1
X_55_ i_pc_change i_reset_n VSS VSS VCC VCC _24_ sky130_fd_sc_hd__or2b_1
X_38_ _06_ i_decode_rs1[3] i_decode_rs1[4] _07_ _08_ VSS VSS VCC VCC _09_
+ sky130_fd_sc_hd__a221o_1
X_54_ inst_sup\[1\] VSS VSS VCC VCC o_inv_inst sky130_fd_sc_hd__inv_2
X_37_ i_alu1_rd[0] i_decode_rs1[0] VSS VSS VCC VCC _08_ sky130_fd_sc_hd__xor2_1
X_53_ _23_ VSS VSS VCC VCC o_decode_stall sky130_fd_sc_hd__inv_2
X_36_ i_alu1_rd[4] VSS VSS VCC VCC _07_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_1_1__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_52_ o_alu1_stall i_need_pause _22_ VSS VSS VCC VCC _23_ sky130_fd_sc_hd__nor3_1
X_35_ i_alu1_rd[3] VSS VSS VCC VCC _06_ sky130_fd_sc_hd__inv_2
X_51_ _12_ _19_ _20_ _02_ _21_ VSS VSS VCC VCC _22_ sky130_fd_sc_hd__a221oi_4
X_34_ _02_ i_decode_rs1[2] i_decode_rs1[1] _04_ VSS VSS VCC VCC _05_ sky130_fd_sc_hd__a2bb2o_1
X_50_ i_alu1_mem_rd VSS VSS VCC VCC _21_ sky130_fd_sc_hd__inv_2
X_33_ i_alu1_rd[1] VSS VSS VCC VCC _04_ sky130_fd_sc_hd__inv_2
X_32_ _02_ i_decode_rs1[2] VSS VSS VCC VCC _03_ sky130_fd_sc_hd__and2_1
X_31_ i_alu1_rd[2] VSS VSS VCC VCC _02_ sky130_fd_sc_hd__inv_2
X_30_ i_alu2_ready VSS VSS VCC VCC o_alu1_stall sky130_fd_sc_hd__clkinv_4
X_69_ o_decode_stall VSS VSS VCC VCC o_fetch_stall sky130_fd_sc_hd__buf_2
X_68_ o_alu2_flush VSS VSS VCC VCC o_decode_flush sky130_fd_sc_hd__buf_2
Xclkbuf_1_0__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_1_0__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_67_ clknet_1_1__leaf_i_clk _01_ VSS VSS VCC VCC inst_sup\[1\] sky130_fd_sc_hd__dfxtp_2
