** sch_path: /media/FlexRV32/asic/blocks/top/top.sch
**.subckt top i_clk i_reset_n
*.ipin i_clk
*.ipin i_reset_n
x1 w_wb_rdata[31] w_wb_rdata[30] w_wb_rdata[29] w_wb_rdata[28] w_wb_rdata[27] w_wb_rdata[26]
+ w_wb_rdata[25] w_wb_rdata[24] w_wb_rdata[23] w_wb_rdata[22] w_wb_rdata[21] w_wb_rdata[20] w_wb_rdata[19]
+ w_wb_rdata[18] w_wb_rdata[17] w_wb_rdata[16] w_wb_rdata[15] w_wb_rdata[14] w_wb_rdata[13] w_wb_rdata[12]
+ w_wb_rdata[11] w_wb_rdata[10] w_wb_rdata[9] w_wb_rdata[8] w_wb_rdata[7] w_wb_rdata[6] w_wb_rdata[5] w_wb_rdata[4]
+ w_wb_rdata[3] w_wb_rdata[2] w_wb_rdata[1] w_wb_rdata[0] w_wb_addr[11] w_wb_addr[10] w_wb_addr[9] w_wb_addr[8]
+ w_wb_addr[7] w_wb_addr[6] w_wb_addr[5] w_wb_addr[4] w_wb_addr[3] w_wb_addr[2] rom
**** begin user architecture code

Xcore_wb VCC VSS i_clk i_reset_n w_wb_we w_wb_sel[0] w_wb_sel[1] w_wb_sel[2] w_wb_sel[3] w_wb_stb
+ w_wb_ack w_wb_cyc  w_wb_addr[0] w_wb_addr[1] w_wb_addr[2] w_wb_addr[3] w_wb_addr[4] w_wb_addr[5]
+ w_wb_addr[6] w_wb_addr[7] w_wb_addr[8] w_wb_addr[9] w_wb_addr[10] w_wb_addr[11] w_wb_addr[12] w_wb_addr[13]
+ w_wb_addr[14] w_wb_addr[15] w_wb_addr[16] w_wb_addr[17] w_wb_addr[18] w_wb_addr[19] w_wb_addr[20] w_wb_addr[21]
+ w_wb_addr[22] w_wb_addr[23] w_wb_addr[24] w_wb_addr[25] w_wb_addr[26] w_wb_addr[27] w_wb_addr[28] w_wb_addr[29]
+ w_wb_addr[30] w_wb_addr[31]  w_wb_wdata[0] w_wb_wdata[1] w_wb_wdata[2] w_wb_wdata[3] w_wb_wdata[4] w_wb_wdata[5]
+ w_wb_wdata[6] w_wb_wdata[7] w_wb_wdata[8] w_wb_wdata[9] w_wb_wdata[10] w_wb_wdata[11] w_wb_wdata[12]
+ w_wb_wdata[13] w_wb_wdata[14] w_wb_wdata[15] w_wb_wdata[16] w_wb_wdata[17] w_wb_wdata[18] w_wb_wdata[19]
+ w_wb_wdata[20] w_wb_wdata[21] w_wb_wdata[22] w_wb_wdata[23] w_wb_wdata[24] w_wb_wdata[25] w_wb_wdata[26]
+ w_wb_wdata[27] w_wb_wdata[28] w_wb_wdata[29] w_wb_wdata[30] w_wb_wdata[31]  w_wb_rdata[0] w_wb_rdata[1]
+ w_wb_rdata[2] w_wb_rdata[3] w_wb_rdata[4] w_wb_rdata[5] w_wb_rdata[6] w_wb_rdata[7] w_wb_rdata[8] w_wb_rdata[9]
+ w_wb_rdata[10] w_wb_rdata[11] w_wb_rdata[12] w_wb_rdata[13] w_wb_rdata[14] w_wb_rdata[15] w_wb_rdata[16]
+ w_wb_rdata[17] w_wb_rdata[18] w_wb_rdata[19] w_wb_rdata[20] w_wb_rdata[21] w_wb_rdata[22] w_wb_rdata[23]
+ w_wb_rdata[24] w_wb_rdata[25] w_wb_rdata[26] w_wb_rdata[27] w_wb_rdata[28] w_wb_rdata[29] w_wb_rdata[30]
+ w_wb_rdata[31]  rv_top_wb

Vw_wb_ack w_wb_ack 0 PWL 0n {VCC}

.include ./rv_top_wb.spice

**** end user architecture code
**.ends

* expanding   symbol:  ../../blocks/rom/rom.sym # of pins=2
** sym_path: /media/FlexRV32/asic/blocks/rom/rom.sym
** sch_path: /media/FlexRV32/asic/blocks/rom/rom.sch
.subckt rom RD[31] RD[30] RD[29] RD[28] RD[27] RD[26] RD[25] RD[24] RD[23] RD[22] RD[21] RD[20]
+ RD[19] RD[18] RD[17] RD[16] RD[15] RD[14] RD[13] RD[12] RD[11] RD[10] RD[9] RD[8] RD[7] RD[6] RD[5] RD[4]
+ RD[3] RD[2] RD[1] RD[0] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0]
*.ipin A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0]
*.opin
*+ RD[31],RD[30],RD[29],RD[28],RD[27],RD[26],RD[25],RD[24],RD[23],RD[22],RD[21],RD[20],RD[19],RD[18],RD[17],RD[16],RD[15],RD[14],RD[13],RD[12],RD[11],RD[10],RD[9],RD[8],RD[7],RD[6],RD[5],RD[4],RD[3],RD[2],RD[1],RD[0]
x1 ROW[255] ROW[254] ROW[253] ROW[252] ROW[251] ROW[250] ROW[249] ROW[248] ROW[247] ROW[246]
+ ROW[245] ROW[244] ROW[243] ROW[242] ROW[241] ROW[240] ROW[239] ROW[238] ROW[237] ROW[236] ROW[235] ROW[234]
+ ROW[233] ROW[232] ROW[231] ROW[230] ROW[229] ROW[228] ROW[227] ROW[226] ROW[225] ROW[224] ROW[223] ROW[222]
+ ROW[221] ROW[220] ROW[219] ROW[218] ROW[217] ROW[216] ROW[215] ROW[214] ROW[213] ROW[212] ROW[211] ROW[210]
+ ROW[209] ROW[208] ROW[207] ROW[206] ROW[205] ROW[204] ROW[203] ROW[202] ROW[201] ROW[200] ROW[199] ROW[198]
+ ROW[197] ROW[196] ROW[195] ROW[194] ROW[193] ROW[192] ROW[191] ROW[190] ROW[189] ROW[188] ROW[187] ROW[186]
+ ROW[185] ROW[184] ROW[183] ROW[182] ROW[181] ROW[180] ROW[179] ROW[178] ROW[177] ROW[176] ROW[175] ROW[174]
+ ROW[173] ROW[172] ROW[171] ROW[170] ROW[169] ROW[168] ROW[167] ROW[166] ROW[165] ROW[164] ROW[163] ROW[162]
+ ROW[161] ROW[160] ROW[159] ROW[158] ROW[157] ROW[156] ROW[155] ROW[154] ROW[153] ROW[152] ROW[151] ROW[150]
+ ROW[149] ROW[148] ROW[147] ROW[146] ROW[145] ROW[144] ROW[143] ROW[142] ROW[141] ROW[140] ROW[139] ROW[138]
+ ROW[137] ROW[136] ROW[135] ROW[134] ROW[133] ROW[132] ROW[131] ROW[130] ROW[129] ROW[128] ROW[127] ROW[126]
+ ROW[125] ROW[124] ROW[123] ROW[122] ROW[121] ROW[120] ROW[119] ROW[118] ROW[117] ROW[116] ROW[115] ROW[114]
+ ROW[113] ROW[112] ROW[111] ROW[110] ROW[109] ROW[108] ROW[107] ROW[106] ROW[105] ROW[104] ROW[103] ROW[102]
+ ROW[101] ROW[100] ROW[99] ROW[98] ROW[97] ROW[96] ROW[95] ROW[94] ROW[93] ROW[92] ROW[91] ROW[90] ROW[89]
+ ROW[88] ROW[87] ROW[86] ROW[85] ROW[84] ROW[83] ROW[82] ROW[81] ROW[80] ROW[79] ROW[78] ROW[77] ROW[76]
+ ROW[75] ROW[74] ROW[73] ROW[72] ROW[71] ROW[70] ROW[69] ROW[68] ROW[67] ROW[66] ROW[65] ROW[64] ROW[63]
+ ROW[62] ROW[61] ROW[60] ROW[59] ROW[58] ROW[57] ROW[56] ROW[55] ROW[54] ROW[53] ROW[52] ROW[51] ROW[50]
+ ROW[49] ROW[48] ROW[47] ROW[46] ROW[45] ROW[44] ROW[43] ROW[42] ROW[41] ROW[40] ROW[39] ROW[38] ROW[37]
+ ROW[36] ROW[35] ROW[34] ROW[33] ROW[32] ROW[31] ROW[30] ROW[29] ROW[28] ROW[27] ROW[26] ROW[25] ROW[24]
+ ROW[23] ROW[22] ROW[21] ROW[20] ROW[19] ROW[18] ROW[17] ROW[16] ROW[15] ROW[14] ROW[13] ROW[12] ROW[11]
+ ROW[10] ROW[9] ROW[8] ROW[7] ROW[6] ROW[5] ROW[4] ROW[3] ROW[2] ROW[1] ROW[0] A[9] A[8] A[7] A[6] A[5] A[4]
+ A[3] A[2] A[1] A[0] COL[3] COL[2] COL[1] COL[0] rom_dec
**** begin user architecture code

.include ../../blocks/rom/rom_data.spice


**** end user architecture code
.ends


* expanding   symbol:  ../../blocks/rom/rom_dec.sym # of pins=3
** sym_path: /media/FlexRV32/asic/blocks/rom/rom_dec.sym
** sch_path: /media/FlexRV32/asic/blocks/rom/rom_dec.sch
.subckt rom_dec ROW[255] ROW[254] ROW[253] ROW[252] ROW[251] ROW[250] ROW[249] ROW[248] ROW[247]
+ ROW[246] ROW[245] ROW[244] ROW[243] ROW[242] ROW[241] ROW[240] ROW[239] ROW[238] ROW[237] ROW[236] ROW[235]
+ ROW[234] ROW[233] ROW[232] ROW[231] ROW[230] ROW[229] ROW[228] ROW[227] ROW[226] ROW[225] ROW[224] ROW[223]
+ ROW[222] ROW[221] ROW[220] ROW[219] ROW[218] ROW[217] ROW[216] ROW[215] ROW[214] ROW[213] ROW[212] ROW[211]
+ ROW[210] ROW[209] ROW[208] ROW[207] ROW[206] ROW[205] ROW[204] ROW[203] ROW[202] ROW[201] ROW[200] ROW[199]
+ ROW[198] ROW[197] ROW[196] ROW[195] ROW[194] ROW[193] ROW[192] ROW[191] ROW[190] ROW[189] ROW[188] ROW[187]
+ ROW[186] ROW[185] ROW[184] ROW[183] ROW[182] ROW[181] ROW[180] ROW[179] ROW[178] ROW[177] ROW[176] ROW[175]
+ ROW[174] ROW[173] ROW[172] ROW[171] ROW[170] ROW[169] ROW[168] ROW[167] ROW[166] ROW[165] ROW[164] ROW[163]
+ ROW[162] ROW[161] ROW[160] ROW[159] ROW[158] ROW[157] ROW[156] ROW[155] ROW[154] ROW[153] ROW[152] ROW[151]
+ ROW[150] ROW[149] ROW[148] ROW[147] ROW[146] ROW[145] ROW[144] ROW[143] ROW[142] ROW[141] ROW[140] ROW[139]
+ ROW[138] ROW[137] ROW[136] ROW[135] ROW[134] ROW[133] ROW[132] ROW[131] ROW[130] ROW[129] ROW[128] ROW[127]
+ ROW[126] ROW[125] ROW[124] ROW[123] ROW[122] ROW[121] ROW[120] ROW[119] ROW[118] ROW[117] ROW[116] ROW[115]
+ ROW[114] ROW[113] ROW[112] ROW[111] ROW[110] ROW[109] ROW[108] ROW[107] ROW[106] ROW[105] ROW[104] ROW[103]
+ ROW[102] ROW[101] ROW[100] ROW[99] ROW[98] ROW[97] ROW[96] ROW[95] ROW[94] ROW[93] ROW[92] ROW[91] ROW[90]
+ ROW[89] ROW[88] ROW[87] ROW[86] ROW[85] ROW[84] ROW[83] ROW[82] ROW[81] ROW[80] ROW[79] ROW[78] ROW[77]
+ ROW[76] ROW[75] ROW[74] ROW[73] ROW[72] ROW[71] ROW[70] ROW[69] ROW[68] ROW[67] ROW[66] ROW[65] ROW[64]
+ ROW[63] ROW[62] ROW[61] ROW[60] ROW[59] ROW[58] ROW[57] ROW[56] ROW[55] ROW[54] ROW[53] ROW[52] ROW[51]
+ ROW[50] ROW[49] ROW[48] ROW[47] ROW[46] ROW[45] ROW[44] ROW[43] ROW[42] ROW[41] ROW[40] ROW[39] ROW[38]
+ ROW[37] ROW[36] ROW[35] ROW[34] ROW[33] ROW[32] ROW[31] ROW[30] ROW[29] ROW[28] ROW[27] ROW[26] ROW[25]
+ ROW[24] ROW[23] ROW[22] ROW[21] ROW[20] ROW[19] ROW[18] ROW[17] ROW[16] ROW[15] ROW[14] ROW[13] ROW[12]
+ ROW[11] ROW[10] ROW[9] ROW[8] ROW[7] ROW[6] ROW[5] ROW[4] ROW[3] ROW[2] ROW[1] ROW[0] A[9] A[8] A[7] A[6]
+ A[5] A[4] A[3] A[2] A[1] A[0] COL[3] COL[2] COL[1] COL[0]
*.ipin A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0]
*.opin
*+ ROW[255],ROW[254],ROW[253],ROW[252],ROW[251],ROW[250],ROW[249],ROW[248],ROW[247],ROW[246],ROW[245],ROW[244],ROW[243],ROW[242],ROW[241],ROW[240],ROW[239],ROW[238],ROW[237],ROW[236],ROW[235],ROW[234],ROW[233],ROW[232],ROW[231],ROW[230],ROW[229],ROW[228],ROW[227],ROW[226],ROW[225],ROW[224],ROW[223],ROW[222],ROW[221],ROW[220],ROW[219],ROW[218],ROW[217],ROW[216],ROW[215],ROW[214],ROW[213],ROW[212],ROW[211],ROW[210],ROW[209],ROW[208],ROW[207],ROW[206],ROW[205],ROW[204],ROW[203],ROW[202],ROW[201],ROW[200],ROW[199],ROW[198],ROW[197],ROW[196],ROW[195],ROW[194],ROW[193],ROW[192],ROW[191],ROW[190],ROW[189],ROW[188],ROW[187],ROW[186],ROW[185],ROW[184],ROW[183],ROW[182],ROW[181],ROW[180],ROW[179],ROW[178],ROW[177],ROW[176],ROW[175],ROW[174],ROW[173],ROW[172],ROW[171],ROW[170],ROW[169],ROW[168],ROW[167],ROW[166],ROW[165],ROW[164],ROW[163],ROW[162],ROW[161],ROW[160],ROW[159],ROW[158],ROW[157],ROW[156],ROW[155],ROW[154],ROW[153],ROW[152],ROW[151],ROW[150],ROW[149],ROW[148],ROW[147],ROW[146],ROW[145],ROW[144],ROW[143],ROW[142],ROW[141],ROW[140],ROW[139],ROW[138],ROW[137],ROW[136],ROW[135],ROW[134],ROW[133],ROW[132],ROW[131],ROW[130],ROW[129],ROW[128],ROW[127],ROW[126],ROW[125],ROW[124],ROW[123],ROW[122],ROW[121],ROW[120],ROW[119],ROW[118],ROW[117],ROW[116],ROW[115],ROW[114],ROW[113],ROW[112],ROW[111],ROW[110],ROW[109],ROW[108],ROW[107],ROW[106],ROW[105],ROW[104],ROW[103],ROW[102],ROW[101],ROW[100],ROW[99],ROW[98],ROW[97],ROW[96],ROW[95],ROW[94],ROW[93],ROW[92],ROW[91],ROW[90],ROW[89],ROW[88],ROW[87],ROW[86],ROW[85],ROW[84],ROW[83],ROW[82],ROW[81],ROW[80],ROW[79],ROW[78],ROW[77],ROW[76],ROW[75],ROW[74],ROW[73],ROW[72],ROW[71],ROW[70],ROW[69],ROW[68],ROW[67],ROW[66],ROW[65],ROW[64],ROW[63],ROW[62],ROW[61],ROW[60],ROW[59],ROW[58],ROW[57],ROW[56],ROW[55],ROW[54],ROW[53],ROW[52],ROW[51],ROW[50],ROW[49],ROW[48],ROW[47],ROW[46],ROW[45],ROW[44],ROW[43],ROW[42],ROW[41],ROW[40],ROW[39],ROW[38],ROW[37],ROW[36],ROW[35],ROW[34],ROW[33],ROW[32],ROW[31],ROW[30],ROW[29],ROW[28],ROW[27],ROW[26],ROW[25],ROW[24],ROW[23],ROW[22],ROW[21],ROW[20],ROW[19],ROW[18],ROW[17],ROW[16],ROW[15],ROW[14],ROW[13],ROW[12],ROW[11],ROW[10],ROW[9],ROW[8],ROW[7],ROW[6],ROW[5],ROW[4],ROW[3],ROW[2],ROW[1],ROW[0]
*.opin COL[3],COL[2],COL[1],COL[0]
x3 net8[1] net8[0] net7[1] net7[0] net9[3] net9[2] net9[1] net9[0] rom_dec_2b
x5 net1[3] net1[2] net1[1] net1[0] ROW[31] ROW[30] ROW[29] ROW[28] ROW[27] ROW[26] ROW[25] ROW[24]
+ ROW[23] ROW[22] ROW[21] ROW[20] ROW[19] ROW[18] ROW[17] ROW[16] SELlo[7] SELlo[6] SELlo[5] SELlo[4]
+ rom_dec_cell
x6 net1[3] net1[2] net1[1] net1[0] ROW[47] ROW[46] ROW[45] ROW[44] ROW[43] ROW[42] ROW[41] ROW[40]
+ ROW[39] ROW[38] ROW[37] ROW[36] ROW[35] ROW[34] ROW[33] ROW[32] SELlo[11] SELlo[10] SELlo[9] SELlo[8]
+ rom_dec_cell
x7 net1[3] net1[2] net1[1] net1[0] ROW[15] ROW[14] ROW[13] ROW[12] ROW[11] ROW[10] ROW[9] ROW[8]
+ ROW[7] ROW[6] ROW[5] ROW[4] ROW[3] ROW[2] ROW[1] ROW[0] SELlo[3] SELlo[2] SELlo[1] SELlo[0] rom_dec_cell
x8 net1[3] net1[2] net1[1] net1[0] ROW[63] ROW[62] ROW[61] ROW[60] ROW[59] ROW[58] ROW[57] ROW[56]
+ ROW[55] ROW[54] ROW[53] ROW[52] ROW[51] ROW[50] ROW[49] ROW[48] SELlo[15] SELlo[14] SELlo[13] SELlo[12]
+ rom_dec_cell
x4 net2[3] net2[2] net2[1] net2[0] ROW[95] ROW[94] ROW[93] ROW[92] ROW[91] ROW[90] ROW[89] ROW[88]
+ ROW[87] ROW[86] ROW[85] ROW[84] ROW[83] ROW[82] ROW[81] ROW[80] SELlo[7] SELlo[6] SELlo[5] SELlo[4]
+ rom_dec_cell
x9 net2[3] net2[2] net2[1] net2[0] ROW[111] ROW[110] ROW[109] ROW[108] ROW[107] ROW[106] ROW[105]
+ ROW[104] ROW[103] ROW[102] ROW[101] ROW[100] ROW[99] ROW[98] ROW[97] ROW[96] SELlo[11] SELlo[10] SELlo[9]
+ SELlo[8] rom_dec_cell
x10 net2[3] net2[2] net2[1] net2[0] ROW[79] ROW[78] ROW[77] ROW[76] ROW[75] ROW[74] ROW[73] ROW[72]
+ ROW[71] ROW[70] ROW[69] ROW[68] ROW[67] ROW[66] ROW[65] ROW[64] SELlo[3] SELlo[2] SELlo[1] SELlo[0]
+ rom_dec_cell
x11 net2[3] net2[2] net2[1] net2[0] ROW[127] ROW[126] ROW[125] ROW[124] ROW[123] ROW[122] ROW[121]
+ ROW[120] ROW[119] ROW[118] ROW[117] ROW[116] ROW[115] ROW[114] ROW[113] ROW[112] SELlo[15] SELlo[14]
+ SELlo[13] SELlo[12] rom_dec_cell
x12 net3[3] net3[2] net3[1] net3[0] ROW[159] ROW[158] ROW[157] ROW[156] ROW[155] ROW[154] ROW[153]
+ ROW[152] ROW[151] ROW[150] ROW[149] ROW[148] ROW[147] ROW[146] ROW[145] ROW[144] SELlo[7] SELlo[6] SELlo[5]
+ SELlo[4] rom_dec_cell
x13 net3[3] net3[2] net3[1] net3[0] ROW[175] ROW[174] ROW[173] ROW[172] ROW[171] ROW[170] ROW[169]
+ ROW[168] ROW[167] ROW[166] ROW[165] ROW[164] ROW[163] ROW[162] ROW[161] ROW[160] SELlo[11] SELlo[10]
+ SELlo[9] SELlo[8] rom_dec_cell
x14 net3[3] net3[2] net3[1] net3[0] ROW[143] ROW[142] ROW[141] ROW[140] ROW[139] ROW[138] ROW[137]
+ ROW[136] ROW[135] ROW[134] ROW[133] ROW[132] ROW[131] ROW[130] ROW[129] ROW[128] SELlo[3] SELlo[2] SELlo[1]
+ SELlo[0] rom_dec_cell
x15 net3[3] net3[2] net3[1] net3[0] ROW[191] ROW[190] ROW[189] ROW[188] ROW[187] ROW[186] ROW[185]
+ ROW[184] ROW[183] ROW[182] ROW[181] ROW[180] ROW[179] ROW[178] ROW[177] ROW[176] SELlo[15] SELlo[14]
+ SELlo[13] SELlo[12] rom_dec_cell
x16 net4[3] net4[2] net4[1] net4[0] ROW[223] ROW[222] ROW[221] ROW[220] ROW[219] ROW[218] ROW[217]
+ ROW[216] ROW[215] ROW[214] ROW[213] ROW[212] ROW[211] ROW[210] ROW[209] ROW[208] SELlo[7] SELlo[6] SELlo[5]
+ SELlo[4] rom_dec_cell
x17 net4[3] net4[2] net4[1] net4[0] ROW[239] ROW[238] ROW[237] ROW[236] ROW[235] ROW[234] ROW[233]
+ ROW[232] ROW[231] ROW[230] ROW[229] ROW[228] ROW[227] ROW[226] ROW[225] ROW[224] SELlo[11] SELlo[10]
+ SELlo[9] SELlo[8] rom_dec_cell
x18 net4[3] net4[2] net4[1] net4[0] ROW[207] ROW[206] ROW[205] ROW[204] ROW[203] ROW[202] ROW[201]
+ ROW[200] ROW[199] ROW[198] ROW[197] ROW[196] ROW[195] ROW[194] ROW[193] ROW[192] SELlo[3] SELlo[2] SELlo[1]
+ SELlo[0] rom_dec_cell
x19 net4[3] net4[2] net4[1] net4[0] ROW[255] ROW[254] ROW[253] ROW[252] ROW[251] ROW[250] ROW[249]
+ ROW[248] ROW[247] ROW[246] ROW[245] ROW[244] ROW[243] ROW[242] ROW[241] ROW[240] SELlo[15] SELlo[14]
+ SELlo[13] SELlo[12] rom_dec_cell
x20 net10[3] net10[2] net10[1] net10[0] SEL_lo[15] SEL_lo[14] SEL_lo[13] SEL_lo[12] SEL_lo[11]
+ SEL_lo[10] SEL_lo[9] SEL_lo[8] SEL_lo[7] SEL_lo[6] SEL_lo[5] SEL_lo[4] SEL_lo[3] SEL_lo[2] SEL_lo[1] SEL_lo[0]
+ net5[3] net5[2] net5[1] net5[0] rom_dec_4b
x21 net11[3] net11[2] net11[1] net11[0] SEL_hi[15] SEL_hi[14] SEL_hi[13] SEL_hi[12] SEL_hi[11]
+ SEL_hi[10] SEL_hi[9] SEL_hi[8] SEL_hi[7] SEL_hi[6] SEL_hi[5] SEL_hi[4] SEL_hi[3] SEL_hi[2] SEL_hi[1] SEL_hi[0]
+ net6[3] net6[2] net6[1] net6[0] rom_dec_4b
x1[1] A[1] VSS VSS VCC VCC net7[1] sky130_fd_sc_hd__inv_8
x1[0] A[0] VSS VSS VCC VCC net7[0] sky130_fd_sc_hd__inv_8
x2[1] net7[1] VSS VSS VCC VCC net8[1] sky130_fd_sc_hd__inv_8
x2[0] net7[0] VSS VSS VCC VCC net8[0] sky130_fd_sc_hd__inv_8
x3[3] net9[3] VSS VSS VCC VCC COL[3] sky130_fd_sc_hd__inv_8
x3[2] net9[2] VSS VSS VCC VCC COL[2] sky130_fd_sc_hd__inv_8
x3[1] net9[1] VSS VSS VCC VCC COL[1] sky130_fd_sc_hd__inv_8
x3[0] net9[0] VSS VSS VCC VCC COL[0] sky130_fd_sc_hd__inv_8
x4[3] A[5] VSS VSS VCC VCC net5[3] sky130_fd_sc_hd__inv_8
x4[2] A[4] VSS VSS VCC VCC net5[2] sky130_fd_sc_hd__inv_8
x4[1] A[3] VSS VSS VCC VCC net5[1] sky130_fd_sc_hd__inv_8
x4[0] A[2] VSS VSS VCC VCC net5[0] sky130_fd_sc_hd__inv_8
x5[3] net5[3] VSS VSS VCC VCC net10[3] sky130_fd_sc_hd__inv_8
x5[2] net5[2] VSS VSS VCC VCC net10[2] sky130_fd_sc_hd__inv_8
x5[1] net5[1] VSS VSS VCC VCC net10[1] sky130_fd_sc_hd__inv_8
x5[0] net5[0] VSS VSS VCC VCC net10[0] sky130_fd_sc_hd__inv_8
x6[3] A[9] VSS VSS VCC VCC net6[3] sky130_fd_sc_hd__inv_8
x6[2] A[8] VSS VSS VCC VCC net6[2] sky130_fd_sc_hd__inv_8
x6[1] A[7] VSS VSS VCC VCC net6[1] sky130_fd_sc_hd__inv_8
x6[0] A[6] VSS VSS VCC VCC net6[0] sky130_fd_sc_hd__inv_8
x7[3] net6[3] VSS VSS VCC VCC net11[3] sky130_fd_sc_hd__inv_8
x7[2] net6[2] VSS VSS VCC VCC net11[2] sky130_fd_sc_hd__inv_8
x7[1] net6[1] VSS VSS VCC VCC net11[1] sky130_fd_sc_hd__inv_8
x7[0] net6[0] VSS VSS VCC VCC net11[0] sky130_fd_sc_hd__inv_8
x18[3] net12[3] VSS VSS VCC VCC SELlo[7] sky130_fd_sc_hd__inv_1
x18[2] net12[2] VSS VSS VCC VCC SELlo[6] sky130_fd_sc_hd__inv_1
x18[1] net12[1] VSS VSS VCC VCC SELlo[5] sky130_fd_sc_hd__inv_1
x18[0] net12[0] VSS VSS VCC VCC SELlo[4] sky130_fd_sc_hd__inv_1
x19[3] net13[3] VSS VSS VCC VCC SELlo[11] sky130_fd_sc_hd__inv_1
x19[2] net13[2] VSS VSS VCC VCC SELlo[10] sky130_fd_sc_hd__inv_1
x19[1] net13[1] VSS VSS VCC VCC SELlo[9] sky130_fd_sc_hd__inv_1
x19[0] net13[0] VSS VSS VCC VCC SELlo[8] sky130_fd_sc_hd__inv_1
x20[3] net14[3] VSS VSS VCC VCC SELlo[15] sky130_fd_sc_hd__inv_1
x20[2] net14[2] VSS VSS VCC VCC SELlo[14] sky130_fd_sc_hd__inv_1
x20[1] net14[1] VSS VSS VCC VCC SELlo[13] sky130_fd_sc_hd__inv_1
x20[0] net14[0] VSS VSS VCC VCC SELlo[12] sky130_fd_sc_hd__inv_1
x21[3] SEL_hi[15] VSS VSS VCC VCC net15[3] sky130_fd_sc_hd__inv_1
x21[2] SEL_hi[14] VSS VSS VCC VCC net15[2] sky130_fd_sc_hd__inv_1
x21[1] SEL_hi[13] VSS VSS VCC VCC net15[1] sky130_fd_sc_hd__inv_1
x21[0] SEL_hi[12] VSS VSS VCC VCC net15[0] sky130_fd_sc_hd__inv_1
x8[3] net15[3] VSS VSS VCC VCC net4[3] sky130_fd_sc_hd__inv_1
x8[2] net15[2] VSS VSS VCC VCC net4[2] sky130_fd_sc_hd__inv_1
x8[1] net15[1] VSS VSS VCC VCC net4[1] sky130_fd_sc_hd__inv_1
x8[0] net15[0] VSS VSS VCC VCC net4[0] sky130_fd_sc_hd__inv_1
x17[3] net16[3] VSS VSS VCC VCC SELlo[3] sky130_fd_sc_hd__inv_4
x17[2] net16[2] VSS VSS VCC VCC SELlo[2] sky130_fd_sc_hd__inv_4
x17[1] net16[1] VSS VSS VCC VCC SELlo[1] sky130_fd_sc_hd__inv_4
x17[0] net16[0] VSS VSS VCC VCC SELlo[0] sky130_fd_sc_hd__inv_4
x22[3] SEL_hi[11] VSS VSS VCC VCC net17[3] sky130_fd_sc_hd__inv_1
x22[2] SEL_hi[10] VSS VSS VCC VCC net17[2] sky130_fd_sc_hd__inv_1
x22[1] SEL_hi[9] VSS VSS VCC VCC net17[1] sky130_fd_sc_hd__inv_1
x22[0] SEL_hi[8] VSS VSS VCC VCC net17[0] sky130_fd_sc_hd__inv_1
x9[3] net17[3] VSS VSS VCC VCC net3[3] sky130_fd_sc_hd__inv_1
x9[2] net17[2] VSS VSS VCC VCC net3[2] sky130_fd_sc_hd__inv_1
x9[1] net17[1] VSS VSS VCC VCC net3[1] sky130_fd_sc_hd__inv_1
x9[0] net17[0] VSS VSS VCC VCC net3[0] sky130_fd_sc_hd__inv_1
x23[3] SEL_hi[7] VSS VSS VCC VCC net18[3] sky130_fd_sc_hd__inv_1
x23[2] SEL_hi[6] VSS VSS VCC VCC net18[2] sky130_fd_sc_hd__inv_1
x23[1] SEL_hi[5] VSS VSS VCC VCC net18[1] sky130_fd_sc_hd__inv_1
x23[0] SEL_hi[4] VSS VSS VCC VCC net18[0] sky130_fd_sc_hd__inv_1
x10[3] net18[3] VSS VSS VCC VCC net2[3] sky130_fd_sc_hd__inv_1
x10[2] net18[2] VSS VSS VCC VCC net2[2] sky130_fd_sc_hd__inv_1
x10[1] net18[1] VSS VSS VCC VCC net2[1] sky130_fd_sc_hd__inv_1
x10[0] net18[0] VSS VSS VCC VCC net2[0] sky130_fd_sc_hd__inv_1
x24[3] SEL_hi[3] VSS VSS VCC VCC net19[3] sky130_fd_sc_hd__inv_1
x24[2] SEL_hi[2] VSS VSS VCC VCC net19[2] sky130_fd_sc_hd__inv_1
x24[1] SEL_hi[1] VSS VSS VCC VCC net19[1] sky130_fd_sc_hd__inv_1
x24[0] SEL_hi[0] VSS VSS VCC VCC net19[0] sky130_fd_sc_hd__inv_1
x11[3] net19[3] VSS VSS VCC VCC net1[3] sky130_fd_sc_hd__inv_4
x11[2] net19[2] VSS VSS VCC VCC net1[2] sky130_fd_sc_hd__inv_4
x11[1] net19[1] VSS VSS VCC VCC net1[1] sky130_fd_sc_hd__inv_4
x11[0] net19[0] VSS VSS VCC VCC net1[0] sky130_fd_sc_hd__inv_4
x13[3] SEL_lo[7] VSS VSS VCC VCC net12[3] sky130_fd_sc_hd__inv_1
x13[2] SEL_lo[6] VSS VSS VCC VCC net12[2] sky130_fd_sc_hd__inv_1
x13[1] SEL_lo[5] VSS VSS VCC VCC net12[1] sky130_fd_sc_hd__inv_1
x13[0] SEL_lo[4] VSS VSS VCC VCC net12[0] sky130_fd_sc_hd__inv_1
x14[3] SEL_lo[11] VSS VSS VCC VCC net13[3] sky130_fd_sc_hd__inv_1
x14[2] SEL_lo[10] VSS VSS VCC VCC net13[2] sky130_fd_sc_hd__inv_1
x14[1] SEL_lo[9] VSS VSS VCC VCC net13[1] sky130_fd_sc_hd__inv_1
x14[0] SEL_lo[8] VSS VSS VCC VCC net13[0] sky130_fd_sc_hd__inv_1
x15[3] SEL_lo[15] VSS VSS VCC VCC net14[3] sky130_fd_sc_hd__inv_1
x15[2] SEL_lo[14] VSS VSS VCC VCC net14[2] sky130_fd_sc_hd__inv_1
x15[1] SEL_lo[13] VSS VSS VCC VCC net14[1] sky130_fd_sc_hd__inv_1
x15[0] SEL_lo[12] VSS VSS VCC VCC net14[0] sky130_fd_sc_hd__inv_1
x12[3] SEL_lo[3] VSS VSS VCC VCC net16[3] sky130_fd_sc_hd__inv_1
x12[2] SEL_lo[2] VSS VSS VCC VCC net16[2] sky130_fd_sc_hd__inv_1
x12[1] SEL_lo[1] VSS VSS VCC VCC net16[1] sky130_fd_sc_hd__inv_1
x12[0] SEL_lo[0] VSS VSS VCC VCC net16[0] sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  ../../blocks/rom/rom_dec_2b.sym # of pins=3
** sym_path: /media/FlexRV32/asic/blocks/rom/rom_dec_2b.sym
** sch_path: /media/FlexRV32/asic/blocks/rom/rom_dec_2b.sch
.subckt rom_dec_2b Ap[1] Ap[0] An[1] An[0] SELn[3] SELn[2] SELn[1] SELn[0]
*.ipin Ap[1],Ap[0]
*.opin SELn[3],SELn[2],SELn[1],SELn[0]
*.ipin An[1],An[0]
x1 An[1] An[0] VSS VSS VCC VCC SELn[0] sky130_fd_sc_hd__nand2_1
x2 An[1] Ap[0] VSS VSS VCC VCC SELn[1] sky130_fd_sc_hd__nand2_1
x3 Ap[1] An[0] VSS VSS VCC VCC SELn[2] sky130_fd_sc_hd__nand2_1
x4 Ap[1] Ap[0] VSS VSS VCC VCC SELn[3] sky130_fd_sc_hd__nand2_1
.ends


* expanding   symbol:  ../../blocks/rom/rom_dec_cell.sym # of pins=3
** sym_path: /media/FlexRV32/asic/blocks/rom/rom_dec_cell.sym
** sch_path: /media/FlexRV32/asic/blocks/rom/rom_dec_cell.sch
.subckt rom_dec_cell ROW[3] ROW[2] ROW[1] ROW[0] SEL[15] SEL[14] SEL[13] SEL[12] SEL[11] SEL[10]
+ SEL[9] SEL[8] SEL[7] SEL[6] SEL[5] SEL[4] SEL[3] SEL[2] SEL[1] SEL[0] COL[3] COL[2] COL[1] COL[0]
*.opin
*+ SEL[15],SEL[14],SEL[13],SEL[12],SEL[11],SEL[10],SEL[9],SEL[8],SEL[7],SEL[6],SEL[5],SEL[4],SEL[3],SEL[2],SEL[1],SEL[0]
*.ipin ROW[3],ROW[2],ROW[1],ROW[0]
*.ipin COL[3],COL[2],COL[1],COL[0]
x2 ROW[1] VSS VSS VCC VCC net3 sky130_fd_sc_hd__inv_2
x3 ROW[2] VSS VSS VCC VCC net2 sky130_fd_sc_hd__inv_2
x4 ROW[3] VSS VSS VCC VCC net1 sky130_fd_sc_hd__inv_2
x5 COL[0] VSS VSS VCC VCC net5 sky130_fd_sc_hd__inv_2
x6 COL[1] VSS VSS VCC VCC net6 sky130_fd_sc_hd__inv_2
x7 COL[2] VSS VSS VCC VCC net7 sky130_fd_sc_hd__inv_2
x8 COL[3] VSS VSS VCC VCC net8 sky130_fd_sc_hd__inv_2
x1 ROW[0] VSS VSS VCC VCC net4 sky130_fd_sc_hd__inv_2
x14 net4 net6 VSS VSS VCC VCC SEL[1] sky130_fd_sc_hd__nand2_1
x15 net3 net6 VSS VSS VCC VCC SEL[5] sky130_fd_sc_hd__nand2_1
x16 net2 net6 VSS VSS VCC VCC SEL[9] sky130_fd_sc_hd__nand2_1
x17 net1 net6 VSS VSS VCC VCC SEL[13] sky130_fd_sc_hd__nand2_1
x18 net4 net5 VSS VSS VCC VCC SEL[0] sky130_fd_sc_hd__nand2_1
x19 net3 net5 VSS VSS VCC VCC SEL[4] sky130_fd_sc_hd__nand2_1
x20 net2 net5 VSS VSS VCC VCC SEL[8] sky130_fd_sc_hd__nand2_1
x21 net1 net5 VSS VSS VCC VCC SEL[12] sky130_fd_sc_hd__nand2_1
x22 net4 net7 VSS VSS VCC VCC SEL[2] sky130_fd_sc_hd__nand2_1
x23 net3 net7 VSS VSS VCC VCC SEL[6] sky130_fd_sc_hd__nand2_1
x24 net2 net7 VSS VSS VCC VCC SEL[10] sky130_fd_sc_hd__nand2_1
x25 net1 net7 VSS VSS VCC VCC SEL[14] sky130_fd_sc_hd__nand2_1
x26 net4 net8 VSS VSS VCC VCC SEL[3] sky130_fd_sc_hd__nand2_1
x27 net3 net8 VSS VSS VCC VCC SEL[7] sky130_fd_sc_hd__nand2_1
x28 net2 net8 VSS VSS VCC VCC SEL[11] sky130_fd_sc_hd__nand2_1
x29 net1 net8 VSS VSS VCC VCC SEL[15] sky130_fd_sc_hd__nand2_1
.ends


* expanding   symbol:  ../../blocks/rom/rom_dec_4b.sym # of pins=3
** sym_path: /media/FlexRV32/asic/blocks/rom/rom_dec_4b.sym
** sch_path: /media/FlexRV32/asic/blocks/rom/rom_dec_4b.sch
.subckt rom_dec_4b Ap[3] Ap[2] Ap[1] Ap[0] SELn[15] SELn[14] SELn[13] SELn[12] SELn[11] SELn[10]
+ SELn[9] SELn[8] SELn[7] SELn[6] SELn[5] SELn[4] SELn[3] SELn[2] SELn[1] SELn[0] An[3] An[2] An[1] An[0]
*.opin
*+ SELn[15],SELn[14],SELn[13],SELn[12],SELn[11],SELn[10],SELn[9],SELn[8],SELn[7],SELn[6],SELn[5],SELn[4],SELn[3],SELn[2],SELn[1],SELn[0]
*.ipin Ap[3],Ap[2],Ap[1],Ap[0]
*.ipin An[3],An[2],An[1],An[0]
x22 An[0] An[1] An[2] An[3] VSS VSS VCC VCC SELn[0] sky130_fd_sc_hd__nand4_1
x23 Ap[0] An[1] An[2] An[3] VSS VSS VCC VCC SELn[1] sky130_fd_sc_hd__nand4_1
x24 An[0] Ap[1] An[2] An[3] VSS VSS VCC VCC SELn[2] sky130_fd_sc_hd__nand4_1
x25 Ap[0] Ap[1] An[2] An[3] VSS VSS VCC VCC SELn[3] sky130_fd_sc_hd__nand4_1
x28 An[0] An[1] Ap[2] An[3] VSS VSS VCC VCC SELn[4] sky130_fd_sc_hd__nand4_1
x29 Ap[0] An[1] Ap[2] An[3] VSS VSS VCC VCC SELn[5] sky130_fd_sc_hd__nand4_1
x30 An[0] Ap[1] Ap[2] An[3] VSS VSS VCC VCC SELn[6] sky130_fd_sc_hd__nand4_1
x31 Ap[0] Ap[1] Ap[2] An[3] VSS VSS VCC VCC SELn[7] sky130_fd_sc_hd__nand4_1
x1 An[0] An[1] An[2] Ap[3] VSS VSS VCC VCC SELn[8] sky130_fd_sc_hd__nand4_1
x2 Ap[0] An[1] An[2] Ap[3] VSS VSS VCC VCC SELn[9] sky130_fd_sc_hd__nand4_1
x3 An[0] Ap[1] An[2] Ap[3] VSS VSS VCC VCC SELn[10] sky130_fd_sc_hd__nand4_1
x4 Ap[0] Ap[1] An[2] Ap[3] VSS VSS VCC VCC SELn[11] sky130_fd_sc_hd__nand4_1
x5 An[0] An[1] Ap[2] Ap[3] VSS VSS VCC VCC SELn[12] sky130_fd_sc_hd__nand4_1
x6 Ap[0] An[1] Ap[2] Ap[3] VSS VSS VCC VCC SELn[13] sky130_fd_sc_hd__nand4_1
x7 An[0] Ap[1] Ap[2] Ap[3] VSS VSS VCC VCC SELn[14] sky130_fd_sc_hd__nand4_1
x8 Ap[0] Ap[1] Ap[2] Ap[3] VSS VSS VCC VCC SELn[15] sky130_fd_sc_hd__nand4_1
.ends

.end
