* NGSPICE file created from rv_alu2.ext - technology: sky130A

.subckt rv_alu2

+ i_clk i_reset_n i_flush
+ i_store i_reg_write i_inst_jal_jalr i_inst_branch i_to_trap
+ i_op1[0] i_op1[1] i_op1[2] i_op1[3] i_op1[4] i_op1[5] i_op1[6] i_op1[7] i_op1[8] i_op1[9] i_op1[10] i_op1[11] i_op1[12] i_op1[13] i_op1[14] i_op1[15] i_op1[16] i_op1[17] i_op1[18] i_op1[19] i_op1[20] i_op1[21] i_op1[22] i_op1[23] i_op1[24] i_op1[25] i_op1[26] i_op1[27] i_op1[28] i_op1[29] i_op1[30] i_op1[31] 
+ i_op2[0] i_op2[1] i_op2[2] i_op2[3] i_op2[4] i_op2[5] i_op2[6] i_op2[7] i_op2[8] i_op2[9] i_op2[10] i_op2[11] i_op2[12] i_op2[13] i_op2[14] i_op2[15] i_op2[16] i_op2[17] i_op2[18] i_op2[19] i_op2[20] i_op2[21] i_op2[22] i_op2[23] i_op2[24] i_op2[25] i_op2[26] i_op2[27] i_op2[28] i_op2[29] i_op2[30] i_op2[31] 
+ i_rd[0] i_rd[1] i_rd[2] i_rd[3] i_rd[4] 
+ i_pc[1] i_pc[2] i_pc[3] i_pc[4] i_pc[5] i_pc[6] i_pc[7] i_pc[8] i_pc[9] i_pc[10] i_pc[11] i_pc[12] i_pc[13] i_pc[14] i_pc[15] 
+ i_pc_next[1] i_pc_next[2] i_pc_next[3] i_pc_next[4] i_pc_next[5] i_pc_next[6] i_pc_next[7] i_pc_next[8] i_pc_next[9] i_pc_next[10] i_pc_next[11] i_pc_next[12] i_pc_next[13] i_pc_next[14] i_pc_next[15] 
+ i_pc_target[1] i_pc_target[2] i_pc_target[3] i_pc_target[4] i_pc_target[5] i_pc_target[6] i_pc_target[7] i_pc_target[8] i_pc_target[9] i_pc_target[10] i_pc_target[11] i_pc_target[12] i_pc_target[13] i_pc_target[14] i_pc_target[15] 
+ i_res_src[0] i_res_src[1] i_res_src[2] 
+ i_funct3[0] i_funct3[1] i_funct3[2] 
+ i_alu_ctrl[0] i_alu_ctrl[1] i_alu_ctrl[2] i_alu_ctrl[3] i_alu_ctrl[4] 
+ i_reg_data2[0] i_reg_data2[1] i_reg_data2[2] i_reg_data2[3] i_reg_data2[4] i_reg_data2[5] i_reg_data2[6] i_reg_data2[7] i_reg_data2[8] i_reg_data2[9] i_reg_data2[10] i_reg_data2[11] i_reg_data2[12] i_reg_data2[13] i_reg_data2[14] i_reg_data2[15] i_reg_data2[16] i_reg_data2[17] i_reg_data2[18] i_reg_data2[19] i_reg_data2[20] i_reg_data2[21] i_reg_data2[22] i_reg_data2[23] i_reg_data2[24] i_reg_data2[25] i_reg_data2[26] i_reg_data2[27] i_reg_data2[28] i_reg_data2[29] i_reg_data2[30] i_reg_data2[31] 
+ i_csr_read
+ i_csr_data[0] i_csr_data[1] i_csr_data[2] i_csr_data[3] i_csr_data[4] i_csr_data[5] i_csr_data[6] i_csr_data[7] i_csr_data[8] i_csr_data[9] i_csr_data[10] i_csr_data[11] i_csr_data[12] i_csr_data[13] i_csr_data[14] i_csr_data[15] i_csr_data[16] i_csr_data[17] i_csr_data[18] i_csr_data[19] i_csr_data[20] i_csr_data[21] i_csr_data[22] i_csr_data[23] i_csr_data[24] i_csr_data[25] i_csr_data[26] i_csr_data[27] i_csr_data[28] i_csr_data[29] i_csr_data[30] i_csr_data[31]
+ o_pc_select o_to_trap
+ o_result[0] o_result[1] o_result[2] o_result[3] o_result[4] o_result[5] o_result[6] o_result[7] o_result[8] o_result[9] o_result[10] o_result[11] o_result[12] o_result[13] o_result[14] o_result[15] o_result[16] o_result[17] o_result[18] o_result[19] o_result[20] o_result[21] o_result[22] o_result[23] o_result[24] o_result[25] o_result[26] o_result[27] o_result[28] o_result[29] o_result[30] o_result[31] 
+ o_add[0] o_add[1] o_add[2] o_add[3] o_add[4] o_add[5] o_add[6] o_add[7] o_add[8] o_add[9] o_add[10] o_add[11] o_add[12] o_add[13] o_add[14] o_add[15] o_add[16] o_add[17] o_add[18] o_add[19] o_add[20] o_add[21] o_add[22] o_add[23] o_add[24] o_add[25] o_add[26] o_add[27] o_add[28] o_add[29] o_add[30] o_add[31]
+ o_store o_reg_write o_ready
+ o_rd[0] o_rd[1] o_rd[2] o_rd[3] o_rd[4] 
+ o_pc_target[1] o_pc_target[2] o_pc_target[3] o_pc_target[4] o_pc_target[5] o_pc_target[6] o_pc_target[7] o_pc_target[8] o_pc_target[9] o_pc_target[10] o_pc_target[11] o_pc_target[12] o_pc_target[13] o_pc_target[14] o_pc_target[15] 
+ o_res_src[2] 
+ o_wdata[0] o_wdata[1] o_wdata[2] o_wdata[3] o_wdata[4] o_wdata[5] o_wdata[6] o_wdata[7] o_wdata[8] o_wdata[9] o_wdata[10] o_wdata[11] o_wdata[12] o_wdata[13] o_wdata[14] o_wdata[15] o_wdata[16] o_wdata[17] o_wdata[18] o_wdata[19] o_wdata[20] o_wdata[21] o_wdata[22] o_wdata[23] o_wdata[24] o_wdata[25] o_wdata[26] o_wdata[27] o_wdata[28] o_wdata[29] o_wdata[30] o_wdata[31]
+ o_data_sel[0] o_wsel[1] o_wsel[2] o_wsel[3] 
+ o_wsel[0] o_funct3[1] o_funct3[2]
+ vccd1 vssd1
X_3155_ _0461_ u_bits.i_op2\[26\] _0465_ u_bits.i_op1\[26\] vssd1 vssd1 vccd1 vccd1
+ _0959_ sky130_fd_sc_hd__a22o_1
X_3086_ _0849_ _0850_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__nand2_1
X_3988_ _1376_ _0909_ _1639_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__mux2_1
X_5727_ clknet_leaf_19_i_clk _0370_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2939_ u_bits.i_op1\[21\] u_bits.i_op1\[22\] _0657_ vssd1 vssd1 vccd1 vccd1 _0752_
+ sky130_fd_sc_hd__mux2_1
X_5658_ clknet_leaf_25_i_clk _0301_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[4\] sky130_fd_sc_hd__dfxtp_1
X_4609_ u_muldiv.divisor\[21\] u_muldiv.dividend\[21\] vssd1 vssd1 vccd1 vccd1 _2032_
+ sky130_fd_sc_hd__or2b_1
X_5589_ clknet_leaf_23_i_clk _0236_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[6\] sky130_fd_sc_hd__dfxtp_1
X_4960_ _2061_ _2065_ _2318_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__a21oi_1
X_4891_ u_muldiv.quotient_msk\[3\] _1210_ _2279_ u_muldiv.quotient_msk\[4\] vssd1
+ vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__a22o_1
X_3911_ _1250_ i_op1[9] _1599_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__mux2_1
X_3842_ _0672_ _1559_ _1560_ _0800_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__o211a_1
X_3773_ _1331_ _1493_ _1495_ _1496_ _0728_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__o221a_1
X_5512_ clknet_leaf_50_i_clk _0160_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[30\]
+ sky130_fd_sc_hd__dfxtp_2
X_2724_ u_muldiv.i_op2_signed alu_ctrl\[2\] vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__or2_2
X_2655_ _0469_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__clkinv_2
X_5443_ clknet_leaf_2_i_clk _0091_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_5374_ clknet_leaf_47_i_clk _0022_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[6\] sky130_fd_sc_hd__dfxtp_1
X_4325_ _1112_ _1847_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__xor2_1
X_4256_ _1802_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_1
X_4187_ _1766_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__clkbuf_1
X_3207_ _0996_ u_bits.i_op2\[27\] _0636_ _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__o22a_1
X_3138_ u_bits.i_op1\[25\] vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__buf_4
X_3069_ _0873_ _0877_ _0524_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_52_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5090_ _2288_ _2437_ vssd1 vssd1 vccd1 vccd1 _2438_ sky130_fd_sc_hd__nor2_1
X_4110_ u_pc_sel.i_pc_next\[15\] i_pc_next[15] _1723_ vssd1 vssd1 vccd1 vccd1 _1728_
+ sky130_fd_sc_hd__mux2_1
X_4041_ _1665_ _1684_ _1685_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__a21o_1
X_4943_ u_muldiv.on_wait vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__clkbuf_4
X_4874_ u_muldiv.quotient_msk\[29\] _2264_ _2229_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__mux2_1
X_3825_ u_bits.i_op2\[17\] _0647_ _0637_ _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__o22a_1
X_3756_ u_muldiv.mul\[44\] _0741_ _1480_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__a21oi_1
X_2707_ _0500_ _0501_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__nand2_1
X_3687_ _1333_ csr_data\[7\] _1388_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__o21ai_1
X_5426_ clknet_leaf_52_i_clk _0074_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[17\] sky130_fd_sc_hd__dfxtp_4
X_2638_ _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__clkbuf_4
X_5357_ clknet_leaf_39_i_clk _0005_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[53\] sky130_fd_sc_hd__dfxtp_1
X_5288_ u_muldiv.divisor\[4\] _2284_ _2285_ u_muldiv.divisor\[5\] vssd1 vssd1 vccd1
+ vccd1 _0395_ sky130_fd_sc_hd__a22o_1
X_4308_ _1831_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__buf_2
X_4239_ _1793_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_1
X_4590_ op_cnt\[0\] op_cnt\[1\] _1204_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__a21oi_1
X_3610_ _1343_ _0861_ _0668_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__mux2_1
X_3541_ u_muldiv.mul\[0\] _0717_ _0719_ u_muldiv.mul\[32\] _1277_ vssd1 vssd1 vccd1
+ vccd1 _1278_ sky130_fd_sc_hd__a221o_1
X_3472_ o_wdata[2] u_wr_mux.i_reg_data2\[18\] _1224_ vssd1 vssd1 vccd1 vccd1 _1227_
+ sky130_fd_sc_hd__mux2_1
X_5211_ _0904_ _2537_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__or2_1
X_5142_ u_muldiv.dividend\[18\] _2484_ _2485_ vssd1 vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__mux2_1
X_5073_ _2422_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__clkbuf_1
X_4024_ _1665_ _1672_ _1673_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__a21o_1
X_4926_ u_muldiv.dividend\[0\] u_muldiv.dividend\[1\] vssd1 vssd1 vccd1 vccd1 _2287_
+ sky130_fd_sc_hd__or2_1
X_4857_ _2161_ _2255_ u_muldiv.o_div\[25\] vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__a21oi_1
X_3808_ _0751_ _1528_ _0712_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__o21a_1
X_4788_ u_muldiv.o_div\[11\] _2194_ u_muldiv.o_div\[12\] vssd1 vssd1 vccd1 vccd1 _2200_
+ sky130_fd_sc_hd__o21ai_1
X_3739_ u_muldiv.dividend\[11\] _1326_ _1327_ u_muldiv.o_div\[11\] _1383_ vssd1 vssd1
+ vccd1 vccd1 _1465_ sky130_fd_sc_hd__a221o_1
X_5409_ clknet_leaf_49_i_clk _0057_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[0\] sky130_fd_sc_hd__dfxtp_1
X_5760_ clknet_leaf_19_i_clk _0403_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_2972_ u_bits.i_op1\[8\] vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__buf_4
X_5691_ clknet_leaf_26_i_clk _0334_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4711_ u_muldiv.divisor\[30\] u_muldiv.dividend\[30\] vssd1 vssd1 vccd1 vccd1 _2134_
+ sky130_fd_sc_hd__xor2_2
X_4642_ _2060_ u_muldiv.dividend\[2\] _2062_ _2063_ _2064_ vssd1 vssd1 vccd1 vccd1
+ _2065_ sky130_fd_sc_hd__a221o_1
X_4573_ o_add[22] _2004_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__and2_1
X_3524_ _0653_ _0647_ _0645_ _0646_ _0650_ _0648_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__mux4_1
X_3455_ u_wr_mux.i_reg_data2\[10\] o_wdata[2] _0718_ vssd1 vssd1 vccd1 vccd1 _1218_
+ sky130_fd_sc_hd__mux2_1
X_3386_ _0523_ _0601_ _0608_ _0612_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__a31o_1
X_5125_ _0647_ _2293_ _2469_ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__nand3_1
X_5056_ _2405_ _2406_ _2375_ vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__a21oi_1
X_4007_ _1641_ _1660_ _1661_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__a21o_1
X_4909_ u_muldiv.quotient_msk\[18\] _2282_ _2281_ u_muldiv.quotient_msk\[19\] vssd1
+ vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__a22o_1
X_3240_ _0747_ _1037_ _1038_ _0453_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__a31o_1
X_3171_ _0825_ _0524_ _0840_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__and3b_1
X_5743_ clknet_leaf_21_i_clk _0386_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[27\]
+ sky130_fd_sc_hd__dfxtp_4
X_2955_ u_bits.i_op1\[21\] vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__buf_4
X_5674_ clknet_leaf_30_i_clk _0317_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[20\] sky130_fd_sc_hd__dfxtp_1
X_2886_ _0698_ _0700_ _0663_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__mux2_1
X_4625_ u_muldiv.divisor\[10\] u_muldiv.dividend\[10\] vssd1 vssd1 vccd1 vccd1 _2048_
+ sky130_fd_sc_hd__or2b_1
X_4556_ _1151_ _2006_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__nor2_1
X_3507_ _1243_ _1245_ vssd1 vssd1 vccd1 vccd1 o_wsel[2] sky130_fd_sc_hd__nor2_4
X_4487_ _1974_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__clkbuf_1
X_3438_ u_muldiv.i_on_end vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__buf_4
X_3369_ _1151_ vssd1 vssd1 vccd1 vccd1 o_add[10] sky130_fd_sc_hd__inv_2
X_5108_ _1878_ _2446_ _2454_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__o21ai_1
X_5039_ u_muldiv.dividend\[9\] _2391_ _2378_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__mux2_1
X_2740_ u_bits.i_op1\[7\] u_muldiv.add_prev\[7\] _0448_ vssd1 vssd1 vccd1 vccd1 _0555_
+ sky130_fd_sc_hd__mux2_1
X_2671_ _0457_ _0485_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__xnor2_1
X_4410_ u_bits.i_op2\[17\] _1915_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__or2_1
X_5390_ clknet_leaf_48_i_clk _0038_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[22\] sky130_fd_sc_hd__dfxtp_2
X_4341_ _0688_ _1859_ _1852_ _1856_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__a31o_1
X_4272_ _1810_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__clkbuf_1
X_3223_ _1021_ _1022_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__and2_1
X_3154_ _0739_ csr_data\[25\] _0958_ _0732_ vssd1 vssd1 vccd1 vccd1 o_result[25] sky130_fd_sc_hd__o211a_2
X_3085_ _0812_ _0853_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__nand2_1
X_3987_ _1641_ _1646_ _1647_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__a21o_1
X_5726_ clknet_leaf_20_i_clk _0369_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_2938_ _0643_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__clkbuf_4
X_5657_ clknet_leaf_25_i_clk _0300_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[3\] sky130_fd_sc_hd__dfxtp_1
X_2869_ _0672_ _0681_ _0683_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__a21oi_1
X_4608_ u_muldiv.divisor\[22\] u_muldiv.dividend\[22\] vssd1 vssd1 vccd1 vccd1 _2031_
+ sky130_fd_sc_hd__and2b_1
X_5588_ clknet_leaf_23_i_clk _0235_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[5\] sky130_fd_sc_hd__dfxtp_1
X_4539_ _2001_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__clkbuf_1
X_4890_ u_muldiv.quotient_msk\[2\] _1210_ _2279_ u_muldiv.quotient_msk\[3\] vssd1
+ vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__a22o_1
X_3910_ _1606_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__clkbuf_1
X_3841_ _0687_ _1318_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__nand2_1
X_3772_ u_muldiv.mul\[13\] _0748_ _1400_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__o21ai_1
X_2723_ _0536_ _0537_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__xor2_4
X_5511_ clknet_leaf_49_i_clk _0159_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[29\]
+ sky130_fd_sc_hd__dfxtp_2
X_2654_ _0467_ _0468_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__xnor2_1
X_5442_ clknet_leaf_1_i_clk _0090_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_5373_ clknet_leaf_47_i_clk _0021_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[5\] sky130_fd_sc_hd__dfxtp_2
X_4324_ _0831_ _1846_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__nand2_1
X_4255_ csr_data\[10\] i_csr_data[10] _1800_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__mux2_1
X_4186_ u_wr_mux.i_reg_data2\[11\] i_reg_data2[11] _1756_ vssd1 vssd1 vccd1 vccd1
+ _1766_ sky130_fd_sc_hd__mux2_1
X_3206_ _0996_ u_bits.i_op2\[27\] _0867_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__a21oi_1
X_3137_ _0644_ _0941_ _0712_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__o21a_1
X_3068_ _0875_ _0876_ _0696_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__mux2_1
X_5709_ clknet_leaf_31_i_clk _0352_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_4040_ u_bits.i_op2\[19\] _1663_ _1675_ i_op2[19] vssd1 vssd1 vccd1 vccd1 _1685_
+ sky130_fd_sc_hd__a22o_1
X_4942_ u_muldiv.dividend\[2\] _2287_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__nand2_1
X_4873_ u_muldiv.o_div\[29\] _1835_ _2264_ _2196_ vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__a31o_1
X_3824_ _0618_ _0639_ _1543_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__and3_1
X_3755_ u_muldiv.dividend\[12\] _0742_ _0743_ u_muldiv.o_div\[12\] _1383_ vssd1 vssd1
+ vccd1 vccd1 _1480_ sky130_fd_sc_hd__a221o_1
X_3686_ _0454_ _1412_ _1414_ _1415_ _1357_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__o221a_1
X_2706_ _0515_ _0519_ _0520_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__o21a_1
X_5425_ clknet_leaf_52_i_clk _0073_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[16\] sky130_fd_sc_hd__dfxtp_4
X_2637_ _0451_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__buf_4
X_5356_ clknet_leaf_39_i_clk _0004_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[52\] sky130_fd_sc_hd__dfxtp_1
X_5287_ u_muldiv.divisor\[3\] _2284_ _2285_ u_muldiv.divisor\[4\] vssd1 vssd1 vccd1
+ vccd1 _0394_ sky130_fd_sc_hd__a22o_1
X_4307_ _1830_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__buf_2
X_4238_ csr_data\[2\] i_csr_data[2] _1789_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__mux2_1
X_4169_ _1757_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__clkbuf_1
X_3540_ u_muldiv.dividend\[0\] _0633_ _0722_ u_muldiv.o_div\[0\] vssd1 vssd1 vccd1
+ vccd1 _1277_ sky130_fd_sc_hd__a22o_1
X_5210_ _2109_ _2546_ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__xnor2_1
X_3471_ _1226_ vssd1 vssd1 vccd1 vccd1 o_wdata[17] sky130_fd_sc_hd__buf_2
X_5141_ _2153_ vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__buf_4
X_5072_ u_muldiv.dividend\[12\] _2421_ _2378_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__mux2_1
X_4023_ u_bits.i_op2\[14\] _1663_ _1651_ i_op2[14] vssd1 vssd1 vccd1 vccd1 _1673_
+ sky130_fd_sc_hd__a22o_1
X_4925_ u_muldiv.dividend\[0\] u_muldiv.dividend\[1\] vssd1 vssd1 vccd1 vccd1 _2286_
+ sky130_fd_sc_hd__nand2_1
X_4856_ u_muldiv.quotient_msk\[25\] _2250_ _2229_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__mux2_1
X_3807_ _0910_ _1262_ _0879_ vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__mux2_1
X_4787_ _2181_ _2197_ _2199_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_51_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3738_ _0714_ _1462_ _1463_ _0623_ _1150_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__o32a_1
X_3669_ _0453_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__clkbuf_2
X_5408_ clknet_leaf_1_i_clk _0056_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_inst_branch
+ sky130_fd_sc_hd__dfxtp_1
X_5339_ _1141_ _1585_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_19_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2971_ _0781_ _0782_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__mux2_2
X_5690_ clknet_leaf_26_i_clk _0333_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4710_ u_muldiv.dividend\[29\] u_muldiv.divisor\[29\] vssd1 vssd1 vccd1 vccd1 _2133_
+ sky130_fd_sc_hd__and2b_1
X_4641_ u_muldiv.divisor\[1\] u_muldiv.dividend\[1\] vssd1 vssd1 vccd1 vccd1 _2064_
+ sky130_fd_sc_hd__and2b_1
X_4572_ _2011_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__clkbuf_1
X_3523_ _1256_ _1259_ _0789_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__mux2_1
X_3454_ _1217_ vssd1 vssd1 vccd1 vccd1 o_wdata[9] sky130_fd_sc_hd__buf_2
X_3385_ _1163_ vssd1 vssd1 vccd1 vccd1 o_add[14] sky130_fd_sc_hd__inv_2
X_5124_ u_bits.i_op1\[15\] u_bits.i_op1\[16\] _2450_ vssd1 vssd1 vccd1 vccd1 _2469_
+ sky130_fd_sc_hd__or3_2
X_5055_ _2047_ _2078_ vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__and2b_1
X_4006_ u_bits.i_op2\[9\] _1637_ _1651_ i_op2[9] vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__a22o_1
X_4908_ u_muldiv.quotient_msk\[17\] _2282_ _2281_ u_muldiv.quotient_msk\[18\] vssd1
+ vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__a22o_1
X_4839_ u_muldiv.o_div\[21\] u_muldiv.o_div\[22\] _2233_ vssd1 vssd1 vccd1 vccd1 _2241_
+ sky130_fd_sc_hd__or3_2
X_3170_ _0836_ _0838_ _0760_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__mux2_1
X_5742_ clknet_leaf_21_i_clk _0385_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[26\]
+ sky130_fd_sc_hd__dfxtp_4
X_2954_ _0751_ _0766_ _0712_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__o21a_1
X_5673_ clknet_leaf_30_i_clk _0316_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[19\] sky130_fd_sc_hd__dfxtp_1
X_2885_ _0699_ u_bits.i_op1\[31\] _0649_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__mux2_1
X_4624_ u_muldiv.dividend\[11\] u_muldiv.divisor\[11\] vssd1 vssd1 vccd1 vccd1 _2047_
+ sky130_fd_sc_hd__and2b_1
X_4555_ _1145_ _2006_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__nor2_1
X_3506_ _1224_ o_add[1] vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__nor2_2
X_4486_ u_muldiv.mul\[3\] u_muldiv.mul\[4\] _1584_ vssd1 vssd1 vccd1 vccd1 _1974_
+ sky130_fd_sc_hd__mux2_1
X_3437_ i_alu_ctrl[1] vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__inv_2
X_3368_ _0589_ _1148_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__xnor2_4
X_5107_ _2303_ _2449_ _2453_ _1829_ vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__a22o_1
X_3299_ _0739_ csr_data\[30\] _1093_ _0732_ vssd1 vssd1 vccd1 vccd1 o_result[30] sky130_fd_sc_hd__o211a_2
X_5038_ _1208_ _2380_ _2381_ _2390_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__a31o_1
X_2670_ _0460_ u_bits.i_op2\[17\] u_bits.i_op1\[17\] _0464_ vssd1 vssd1 vccd1 vccd1
+ _0485_ sky130_fd_sc_hd__a22o_1
X_4340_ _1859_ _1850_ _0688_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__a21oi_1
X_4271_ csr_data\[18\] i_csr_data[18] _1800_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__mux2_1
X_3222_ _1019_ _1020_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__or2_1
X_3153_ _0939_ _0957_ _0447_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__a21o_1
X_3084_ u_muldiv.mul\[24\] _0740_ _0741_ u_muldiv.mul\[56\] _0891_ vssd1 vssd1 vccd1
+ vccd1 _0892_ sky130_fd_sc_hd__a221o_1
X_3986_ _0909_ _1637_ _1638_ i_op2[3] vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__a22o_1
X_5725_ clknet_leaf_26_i_clk _0368_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2937_ _0749_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__buf_2
X_5656_ clknet_leaf_24_i_clk _0299_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[2\] sky130_fd_sc_hd__dfxtp_1
X_4607_ u_muldiv.divisor\[28\] u_muldiv.dividend\[28\] vssd1 vssd1 vccd1 vccd1 _2030_
+ sky130_fd_sc_hd__nand2b_4
X_2868_ _0625_ _0682_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__nand2_1
X_5587_ clknet_leaf_23_i_clk _0234_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[4\] sky130_fd_sc_hd__dfxtp_1
X_2799_ _0523_ _0601_ _0608_ _0613_ _0484_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__a311o_1
X_4538_ u_muldiv.mul\[28\] u_muldiv.mul\[29\] _1583_ vssd1 vssd1 vccd1 vccd1 _2001_
+ sky130_fd_sc_hd__mux2_1
X_4469_ u_bits.i_op2\[29\] _1852_ _1962_ _1831_ vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__a31o_1
X_3840_ _0833_ _0835_ _0836_ _0838_ _0825_ _0707_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__mux4_1
X_3771_ u_muldiv.mul\[45\] _0741_ _1494_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__a21oi_1
X_2722_ u_bits.i_op1\[1\] u_muldiv.add_prev\[1\] _0449_ vssd1 vssd1 vccd1 vccd1 _0537_
+ sky130_fd_sc_hd__mux2_2
X_5510_ clknet_leaf_49_i_clk _0158_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[28\]
+ sky130_fd_sc_hd__dfxtp_2
X_2653_ u_bits.i_op1\[20\] u_muldiv.add_prev\[20\] _0451_ vssd1 vssd1 vccd1 vccd1
+ _0468_ sky130_fd_sc_hd__mux2_1
X_5441_ clknet_leaf_1_i_clk _0089_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_5372_ clknet_leaf_47_i_clk _0020_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[4\] sky130_fd_sc_hd__dfxtp_2
X_4323_ _1845_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__buf_2
X_4254_ _1801_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
X_4185_ _1765_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__clkbuf_1
X_3205_ _0674_ _1004_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__a21o_1
X_3136_ _0909_ _0940_ _0911_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__o21a_1
X_3067_ u_bits.i_op1\[11\] u_bits.i_op1\[10\] u_bits.i_op1\[9\] u_bits.i_op1\[8\]
+ _0657_ _0663_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__mux4_1
X_5708_ clknet_leaf_30_i_clk _0351_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_3969_ i_rd[3] _1632_ _1636_ o_rd[3] vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__a22o_1
X_5639_ clknet_leaf_41_i_clk _0286_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_4941_ u_muldiv.dividend\[0\] u_muldiv.dividend\[1\] u_muldiv.dividend\[2\] vssd1
+ vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__or3_1
X_4872_ _2267_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__clkbuf_1
X_3823_ u_bits.i_op2\[17\] _0647_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__nand2_1
X_3754_ _0714_ _1477_ _1478_ _0623_ _1157_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__o32a_1
X_3685_ u_muldiv.mul\[7\] _1330_ _1400_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__o21ai_1
X_2705_ _0513_ _0514_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__nand2_1
X_2636_ _0450_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__clkbuf_4
X_5424_ clknet_leaf_52_i_clk _0072_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[15\] sky130_fd_sc_hd__dfxtp_4
X_5355_ _0616_ _2004_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__nor2_1
X_5286_ u_muldiv.divisor\[2\] _2284_ _2285_ u_muldiv.divisor\[3\] vssd1 vssd1 vccd1
+ vccd1 _0393_ sky130_fd_sc_hd__a22o_1
X_4306_ u_muldiv.on_wait u_muldiv.i_on_end vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__or2_1
X_4237_ _1792_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__clkbuf_1
X_4168_ o_wdata[2] i_reg_data2[2] _1756_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__mux2_1
X_4099_ u_pc_sel.i_pc_next\[10\] i_pc_next[10] _1712_ vssd1 vssd1 vccd1 vccd1 _1722_
+ sky130_fd_sc_hd__mux2_1
X_3119_ _0636_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__clkbuf_4
X_3470_ o_wdata[1] u_wr_mux.i_reg_data2\[17\] _1224_ vssd1 vssd1 vccd1 vccd1 _1226_
+ sky130_fd_sc_hd__mux2_1
X_5140_ _2476_ _2483_ _1877_ vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__mux2_1
X_5071_ _2414_ _2420_ _1877_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__mux2_1
X_4022_ u_bits.i_op2\[15\] _1487_ _1657_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__mux2_1
X_4924_ u_muldiv.quotient_msk\[30\] _2284_ _2285_ u_muldiv.quotient_msk\[31\] vssd1
+ vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__a22o_1
X_4855_ u_muldiv.o_div\[25\] _2170_ _2250_ _2196_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__a31o_1
X_4786_ _2167_ _2198_ u_muldiv.o_div\[11\] vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__a21oi_1
X_3806_ u_muldiv.mul\[16\] _0717_ _0720_ u_muldiv.mul\[48\] _1526_ vssd1 vssd1 vccd1
+ vccd1 _1527_ sky130_fd_sc_hd__a221o_1
X_3737_ u_bits.i_op2\[11\] _1251_ _0906_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__a21oi_1
X_3668_ u_muldiv.mul\[38\] _1325_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__a21oi_1
X_3599_ _0454_ _1324_ _1329_ _1332_ _1333_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__o221a_1
X_5407_ clknet_leaf_1_i_clk _0055_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_inst_jal_jalr
+ sky130_fd_sc_hd__dfxtp_1
X_5338_ _1142_ _1585_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__nor2_1
X_5269_ u_muldiv.dividend\[30\] _2583_ vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__nor2_1
X_2970_ _0663_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__clkbuf_4
X_4640_ u_muldiv.dividend\[0\] u_muldiv.divisor\[0\] vssd1 vssd1 vccd1 vccd1 _2063_
+ sky130_fd_sc_hd__or2b_1
X_4571_ o_add[21] _2004_ vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__and2_1
X_3522_ u_bits.i_op1\[4\] _1257_ _0786_ _1258_ _0651_ _0783_ vssd1 vssd1 vccd1 vccd1
+ _1259_ sky130_fd_sc_hd__mux4_1
X_3453_ u_wr_mux.i_reg_data2\[9\] o_wdata[1] _0718_ vssd1 vssd1 vccd1 vccd1 _1217_
+ sky130_fd_sc_hd__mux2_1
X_5123_ u_muldiv.dividend\[17\] u_muldiv.dividend\[16\] _2444_ vssd1 vssd1 vccd1 vccd1
+ _2468_ sky130_fd_sc_hd__or3_2
X_3384_ _0509_ _1160_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__xor2_4
X_5054_ _2048_ _2397_ vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__and2_1
X_4005_ _1445_ u_bits.i_op2\[8\] _1657_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__mux2_1
X_4907_ _1209_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__buf_2
X_4838_ u_muldiv.o_div\[21\] _2233_ u_muldiv.o_div\[22\] vssd1 vssd1 vccd1 vccd1 _2240_
+ sky130_fd_sc_hd__o21ai_1
X_4769_ u_muldiv.o_div\[7\] _2179_ u_muldiv.o_div\[8\] vssd1 vssd1 vccd1 vccd1 _2185_
+ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_50_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5741_ clknet_leaf_21_i_clk _0384_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[25\]
+ sky130_fd_sc_hd__dfxtp_2
X_2953_ _0759_ _0765_ _0707_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__mux2_1
X_5672_ clknet_leaf_28_i_clk _0315_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[18\] sky130_fd_sc_hd__dfxtp_1
X_2884_ u_bits.i_op1\[30\] vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__clkbuf_4
X_4623_ _2044_ _2045_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__nand2_1
X_4554_ _1147_ _2006_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__nor2_1
X_3505_ _1242_ _1244_ vssd1 vssd1 vccd1 vccd1 o_wsel[1] sky130_fd_sc_hd__nor2_4
X_4485_ _1973_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_1
X_3436_ _1204_ _1192_ _1203_ vssd1 vssd1 vccd1 vccd1 mul_op2_signed_next sky130_fd_sc_hd__nor3_1
X_3367_ _1150_ vssd1 vssd1 vccd1 vccd1 o_add[11] sky130_fd_sc_hd__inv_2
X_5106_ _1206_ _2451_ _2452_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__or3_1
X_5037_ _2303_ _2384_ _2389_ vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__a21oi_1
X_3298_ _1079_ _1092_ _0446_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_18_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4270_ _1809_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__clkbuf_1
X_3221_ _1019_ _1020_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__nand2_1
X_3152_ _0750_ o_add[25] _0954_ _0956_ _0804_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__a221o_1
X_3083_ u_muldiv.dividend\[24\] _0742_ _0743_ u_muldiv.o_div\[24\] _0744_ vssd1 vssd1
+ vccd1 vccd1 _0891_ sky130_fd_sc_hd__a221o_1
X_3985_ _0688_ _0923_ _1639_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__mux2_1
X_5724_ clknet_leaf_26_i_clk _0367_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_2936_ _0747_ _0748_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__nand2_2
X_5655_ clknet_leaf_31_i_clk _0298_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[1\] sky130_fd_sc_hd__dfxtp_1
X_2867_ o_funct3[1] o_funct3[0] vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__and2b_1
X_4606_ _1835_ _2026_ _2027_ _2028_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__a31o_1
X_5586_ clknet_leaf_23_i_clk _0233_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[3\] sky130_fd_sc_hd__dfxtp_1
X_2798_ _0610_ _0612_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__or2_1
X_4537_ _2000_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__clkbuf_1
X_4468_ _1850_ _1962_ u_bits.i_op2\[29\] vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__a21oi_1
X_3419_ _1171_ _1188_ _0618_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__a21oi_1
X_4399_ u_bits.i_op2\[15\] _1852_ _1906_ _1856_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__a31o_1
X_3770_ u_muldiv.dividend\[13\] _0742_ _0743_ u_muldiv.o_div\[13\] _1383_ vssd1 vssd1
+ vccd1 vccd1 _1494_ sky130_fd_sc_hd__a221o_1
X_2721_ _0456_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__xnor2_2
X_5440_ clknet_leaf_0_i_clk _0088_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[31\] sky130_fd_sc_hd__dfxtp_4
X_2652_ _0458_ _0466_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__xnor2_2
X_5371_ clknet_leaf_46_i_clk _0019_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[3\] sky130_fd_sc_hd__dfxtp_2
X_4322_ _1844_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__buf_2
X_4253_ csr_data\[9\] i_csr_data[9] _1800_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__mux2_1
X_3204_ _0669_ _0788_ _0881_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__and3b_1
X_4184_ u_wr_mux.i_reg_data2\[10\] i_reg_data2[10] _1756_ vssd1 vssd1 vccd1 vccd1
+ _1765_ sky130_fd_sc_hd__mux2_1
X_3135_ _0757_ _0764_ _0696_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__mux2_1
X_3066_ _0782_ _0874_ _0533_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__mux2_1
X_3968_ i_rd[2] _1632_ _1636_ o_rd[2] vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__a22o_1
X_5707_ clknet_leaf_30_i_clk _0350_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_2919_ _0461_ u_bits.i_op2\[21\] _0465_ u_bits.i_op1\[21\] vssd1 vssd1 vccd1 vccd1
+ _0733_ sky130_fd_sc_hd__a22o_1
X_3899_ _0794_ i_op1[3] _1599_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__mux2_1
X_5638_ clknet_leaf_41_i_clk _0285_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_5569_ clknet_leaf_9_i_clk _0216_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_4940_ _2300_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__clkbuf_1
X_4871_ u_muldiv.o_div\[28\] _2266_ _2244_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__mux2_1
X_3822_ _0751_ _1290_ _0711_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__o21a_1
X_3753_ u_bits.i_op2\[12\] _0777_ _0906_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__a21oi_1
X_3684_ u_muldiv.mul\[39\] _1325_ _1413_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__a21oi_1
X_2704_ _0517_ _0518_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__nand2_1
X_2635_ _0449_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__buf_4
X_5423_ clknet_leaf_52_i_clk _0071_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[14\] sky130_fd_sc_hd__dfxtp_4
X_5354_ _2630_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__clkbuf_1
X_4305_ _1828_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__clkbuf_4
X_5285_ u_muldiv.divisor\[1\] _2284_ _2285_ u_muldiv.divisor\[2\] vssd1 vssd1 vccd1
+ vccd1 _0392_ sky130_fd_sc_hd__a22o_1
X_4236_ csr_data\[1\] i_csr_data[1] _1789_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__mux2_1
X_4167_ _1711_ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__clkbuf_4
X_3118_ _0642_ _0683_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__nor2_4
X_4098_ _1721_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__clkbuf_1
X_3049_ _0627_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__buf_2
X_5070_ _1826_ _2415_ _2416_ _2418_ _2419_ vssd1 vssd1 vccd1 vccd1 _2420_ sky130_fd_sc_hd__a32o_1
X_4021_ _1665_ _1670_ _1671_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__a21o_1
X_4923_ _1946_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__clkbuf_4
X_4854_ _2253_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__clkbuf_1
X_4785_ u_muldiv.quotient_msk\[11\] _2194_ _2156_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__mux2_1
X_3805_ u_muldiv.dividend\[16\] _0721_ _0723_ u_muldiv.o_div\[16\] _0724_ vssd1 vssd1
+ vccd1 vccd1 _1526_ sky130_fd_sc_hd__a221o_1
X_3736_ _0908_ _1461_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__nor2_1
X_3667_ u_muldiv.dividend\[6\] _1326_ _1327_ u_muldiv.o_div\[6\] _1383_ vssd1 vssd1
+ vccd1 vccd1 _1398_ sky130_fd_sc_hd__a221o_1
X_3598_ _0728_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__buf_2
X_5406_ clknet_leaf_51_i_clk _0054_ vssd1 vssd1 vccd1 vccd1 o_rd[4] sky130_fd_sc_hd__dfxtp_2
X_5337_ _1135_ _1585_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__nor2_1
X_5268_ _2375_ _2595_ _2596_ _2597_ _2599_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__a32o_1
X_4219_ _1783_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__clkbuf_1
X_5199_ u_bits.i_op1\[21\] _0691_ _0692_ _2511_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__or4_2
X_4570_ _0616_ _2007_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__nor2_1
X_3521_ u_bits.i_op1\[7\] vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__clkbuf_4
X_3452_ _1216_ vssd1 vssd1 vccd1 vccd1 o_wdata[8] sky130_fd_sc_hd__buf_2
X_3383_ _1162_ vssd1 vssd1 vccd1 vccd1 o_add[15] sky130_fd_sc_hd__inv_2
X_5122_ u_muldiv.dividend\[16\] _2444_ u_muldiv.dividend\[17\] vssd1 vssd1 vccd1 vccd1
+ _2467_ sky130_fd_sc_hd__o21ai_1
X_5053_ u_muldiv.dividend\[10\] _2380_ u_muldiv.dividend\[11\] vssd1 vssd1 vccd1 vccd1
+ _2404_ sky130_fd_sc_hd__o21ai_1
X_4004_ _1641_ _1658_ _1659_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__a21o_1
X_4906_ u_muldiv.quotient_msk\[16\] _2280_ _2281_ u_muldiv.quotient_msk\[17\] vssd1
+ vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__a22o_1
X_4837_ _2181_ _2237_ _2239_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__a21oi_1
X_4768_ _2181_ _2182_ _2184_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__a21oi_1
X_4699_ _2031_ _2105_ _2106_ _2119_ _2121_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__o311a_1
X_3719_ _1445_ _1305_ _1267_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__a21oi_1
X_5740_ clknet_leaf_17_i_clk _0383_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[24\]
+ sky130_fd_sc_hd__dfxtp_4
X_2952_ _0760_ _0764_ _0704_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__o21a_1
X_5671_ clknet_leaf_31_i_clk _0314_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[17\] sky130_fd_sc_hd__dfxtp_1
X_2883_ u_bits.i_op1\[28\] _0697_ _0649_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__mux2_1
X_4622_ u_muldiv.dividend\[12\] u_muldiv.divisor\[12\] vssd1 vssd1 vccd1 vccd1 _2045_
+ sky130_fd_sc_hd__or2b_1
X_4553_ _1141_ _2006_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__nor2_1
X_4484_ u_muldiv.mul\[2\] u_muldiv.mul\[3\] _1584_ vssd1 vssd1 vccd1 vccd1 _1973_
+ sky130_fd_sc_hd__mux2_1
X_3504_ _0621_ o_add[0] vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__nor2_2
X_3435_ o_ready vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__clkbuf_4
X_3366_ _0584_ _1149_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__xnor2_4
X_5105_ _2293_ _2450_ _0654_ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__a21oi_1
X_3297_ _0750_ o_add[30] _1090_ _1091_ _0804_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__a221o_1
X_5036_ _1206_ _2387_ _2388_ _1828_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__o31a_1
X_3220_ u_bits.i_op1\[28\] u_muldiv.add_prev\[28\] _0452_ vssd1 vssd1 vccd1 vccd1
+ _1020_ sky130_fd_sc_hd__mux2_1
X_3151_ _0629_ _0950_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__a21oi_1
X_3082_ _0739_ csr_data\[23\] _0890_ vssd1 vssd1 vccd1 vccd1 o_result[23] sky130_fd_sc_hd__o21a_2
X_3984_ _1641_ _1644_ _1645_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__a21o_1
X_5723_ clknet_leaf_26_i_clk _0366_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2935_ _0625_ _0639_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__nand2_2
X_5654_ clknet_leaf_22_i_clk u_muldiv.i_on_wait vssd1 vssd1 vccd1 vccd1 u_muldiv.on_wait
+ sky130_fd_sc_hd__dfxtp_2
X_2866_ _0674_ _0680_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__nand2_1
X_4605_ u_muldiv.quotient_msk\[1\] u_muldiv.o_div\[1\] _1841_ vssd1 vssd1 vccd1 vccd1
+ _2028_ sky130_fd_sc_hd__o21a_1
X_5585_ clknet_leaf_23_i_clk _0232_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[2\] sky130_fd_sc_hd__dfxtp_1
X_2797_ _0492_ _0611_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__nand2_2
X_4536_ u_muldiv.mul\[27\] u_muldiv.mul\[28\] _1989_ vssd1 vssd1 vccd1 vccd1 _2000_
+ sky130_fd_sc_hd__mux2_1
X_4467_ u_bits.i_op2\[28\] _1958_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__or2_1
X_4398_ _1868_ _1906_ u_bits.i_op2\[15\] vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__a21oi_1
X_3418_ _1171_ _1188_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__or2_1
X_3349_ _1137_ vssd1 vssd1 vccd1 vccd1 o_add[4] sky130_fd_sc_hd__inv_2
X_5019_ _1258_ _2363_ _2293_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__o21ai_1
X_2720_ _0448_ u_bits.i_op1\[1\] _0497_ _0534_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__a31o_1
X_2651_ _0461_ u_bits.i_op2\[20\] _0465_ u_bits.i_op1\[20\] vssd1 vssd1 vccd1 vccd1
+ _0466_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_17_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5370_ clknet_leaf_47_i_clk _0018_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[2\] sky130_fd_sc_hd__dfxtp_2
X_4321_ _0620_ u_bits.i_op2\[31\] vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__and2b_1
X_4252_ _1711_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__clkbuf_4
X_3203_ _0876_ _0880_ _0825_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__mux2_1
X_4183_ _1764_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__clkbuf_1
X_3134_ u_muldiv.mul\[25\] _0740_ _0741_ u_muldiv.mul\[57\] _0938_ vssd1 vssd1 vccd1
+ vccd1 _0939_ sky130_fd_sc_hd__a221o_1
X_3065_ u_bits.i_op1\[13\] u_bits.i_op1\[12\] _0656_ vssd1 vssd1 vccd1 vccd1 _0874_
+ sky130_fd_sc_hd__mux2_1
X_3967_ i_rd[1] _1632_ _1636_ o_rd[1] vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__a22o_1
X_5706_ clknet_leaf_30_i_clk _0349_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_2918_ _0447_ _0727_ _0729_ _0732_ vssd1 vssd1 vccd1 vccd1 o_result[20] sky130_fd_sc_hd__o211a_2
X_3898_ _1600_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__clkbuf_1
X_2849_ _0661_ _0662_ _0663_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__mux2_1
X_5637_ clknet_leaf_41_i_clk _0284_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_5568_ clknet_leaf_3_i_clk _0215_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_4519_ _1991_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__clkbuf_1
X_5499_ clknet_leaf_43_i_clk _0147_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_4870_ _2208_ _2263_ _2264_ _2265_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__a31o_1
X_3821_ u_muldiv.mul\[17\] _0717_ _0720_ u_muldiv.mul\[49\] _1540_ vssd1 vssd1 vccd1
+ vccd1 _1541_ sky130_fd_sc_hd__a221o_1
X_3752_ _0908_ _1476_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__nor2_1
X_3683_ u_muldiv.dividend\[7\] _1326_ _1327_ u_muldiv.o_div\[7\] _1383_ vssd1 vssd1
+ vccd1 vccd1 _1413_ sky130_fd_sc_hd__a221o_1
X_2703_ u_bits.i_op1\[12\] u_muldiv.add_prev\[12\] _0450_ vssd1 vssd1 vccd1 vccd1
+ _0518_ sky130_fd_sc_hd__mux2_1
X_2634_ _0448_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__clkbuf_4
X_5422_ clknet_leaf_48_i_clk _0070_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[13\] sky130_fd_sc_hd__dfxtp_1
X_5353_ o_add[19] _1214_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__and2_1
X_4304_ _1826_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__nand2_2
X_5284_ u_muldiv.divisor\[0\] _2284_ _2285_ u_muldiv.divisor\[1\] vssd1 vssd1 vccd1
+ vccd1 _0391_ sky130_fd_sc_hd__a22o_1
X_4235_ _1791_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__clkbuf_1
X_4166_ _1755_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__clkbuf_1
X_3117_ _0660_ _0922_ _0664_ _0652_ _0879_ _0923_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__mux4_1
X_4097_ u_pc_sel.i_pc_next\[9\] i_pc_next[9] _1712_ vssd1 vssd1 vccd1 vccd1 _1721_
+ sky130_fd_sc_hd__mux2_1
X_3048_ u_muldiv.mul\[23\] _0717_ _0720_ u_muldiv.mul\[55\] _0856_ vssd1 vssd1 vccd1
+ vccd1 _0857_ sky130_fd_sc_hd__a221o_1
X_4999_ u_muldiv.dividend\[6\] _2354_ _2244_ vssd1 vssd1 vccd1 vccd1 _2355_ sky130_fd_sc_hd__mux2_1
X_4020_ _1487_ _1663_ _1651_ i_op2[13] vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__a22o_1
X_4922_ u_muldiv.quotient_msk\[29\] _2284_ _2283_ u_muldiv.quotient_msk\[30\] vssd1
+ vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__a22o_1
X_4853_ u_muldiv.o_div\[24\] _2252_ _2244_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__mux2_1
X_4784_ _2170_ u_muldiv.o_div\[11\] _2194_ _2196_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__a31o_1
X_3804_ _1524_ _1525_ _0730_ u_pc_sel.i_pc_next\[15\] vssd1 vssd1 vccd1 vccd1 o_result[15]
+ sky130_fd_sc_hd__a2bb2o_2
X_3735_ _1110_ _1006_ _1458_ _1248_ _1460_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__a221o_1
X_5405_ clknet_leaf_51_i_clk _0053_ vssd1 vssd1 vccd1 vccd1 o_rd[3] sky130_fd_sc_hd__dfxtp_2
X_3666_ _1274_ _1395_ _1396_ _0624_ _1142_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__o32a_1
X_3597_ u_muldiv.mul\[2\] _1330_ _1331_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__o21ai_1
X_5336_ _1137_ _1585_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__nor2_1
X_5267_ _2134_ _2598_ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__nand2_1
X_4218_ u_wr_mux.i_reg_data2\[26\] i_reg_data2[26] _1778_ vssd1 vssd1 vccd1 vccd1
+ _1783_ sky130_fd_sc_hd__mux2_1
X_5198_ u_muldiv.dividend\[24\] _2525_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__xor2_1
X_4149_ _1224_ i_funct3[1] _1745_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__mux2_1
X_3520_ u_bits.i_op1\[5\] vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__clkbuf_4
X_3451_ u_wr_mux.i_reg_data2\[8\] o_wdata[0] _0718_ vssd1 vssd1 vccd1 vccd1 _1216_
+ sky130_fd_sc_hd__mux2_1
X_3382_ _1158_ _1161_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__xor2_4
X_5121_ _2092_ _2465_ vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__xnor2_1
X_5052_ u_muldiv.dividend\[11\] u_muldiv.dividend\[10\] _2380_ vssd1 vssd1 vccd1 vccd1
+ _2403_ sky130_fd_sc_hd__or3_2
X_4003_ u_bits.i_op2\[8\] _1637_ _1651_ i_op2[8] vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__a22o_1
X_4905_ u_muldiv.quotient_msk\[15\] _2280_ _2281_ u_muldiv.quotient_msk\[16\] vssd1
+ vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__a22o_1
X_4836_ _2161_ _2238_ u_muldiv.o_div\[21\] vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__a21oi_1
X_4767_ _2167_ _2183_ u_muldiv.o_div\[7\] vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__a21oi_1
X_4698_ _2120_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__inv_2
X_3718_ u_bits.i_op2\[10\] vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__clkbuf_4
X_3649_ _1376_ _1257_ _1272_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__a21oi_1
X_5319_ _0702_ _1969_ u_bits.i_op2\[31\] vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__a21o_1
X_2951_ _0659_ _0761_ _0762_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__o22a_1
X_5670_ clknet_leaf_30_i_clk _0313_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[16\] sky130_fd_sc_hd__dfxtp_1
X_4621_ u_muldiv.divisor\[12\] u_muldiv.dividend\[12\] vssd1 vssd1 vccd1 vccd1 _2044_
+ sky130_fd_sc_hd__or2b_1
X_2882_ u_bits.i_op1\[29\] vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__buf_4
X_4552_ _1142_ _2006_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__nor2_1
X_4483_ _1972_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_1
X_3503_ _1242_ _1243_ vssd1 vssd1 vccd1 vccd1 o_wsel[0] sky130_fd_sc_hd__nor2_4
X_3434_ i_flush _1203_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__nor2_1
X_3365_ _0589_ _1148_ _0603_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__a21bo_1
X_5104_ _0654_ _2292_ _2450_ vssd1 vssd1 vccd1 vccd1 _2451_ sky130_fd_sc_hd__and3_1
X_3296_ _0629_ _1086_ _0955_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__a21oi_1
X_5035_ _2295_ _2386_ _1250_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__a21oi_1
X_4819_ u_muldiv.o_div\[17\] _2218_ u_muldiv.o_div\[18\] vssd1 vssd1 vccd1 vccd1 _2225_
+ sky130_fd_sc_hd__o21ai_1
X_5799_ clknet_leaf_34_i_clk _0441_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[47\] sky130_fd_sc_hd__dfxtp_1
X_3150_ u_mux.i_add_override vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__buf_2
X_3081_ _0730_ _0889_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__nor2_1
X_5722_ clknet_leaf_25_i_clk _0365_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3983_ _0923_ _1637_ _1638_ i_op2[2] vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__a22o_1
X_2934_ u_mux.i_add_override vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__clkinv_2
X_5653_ clknet_leaf_10_i_clk _0297_ vssd1 vssd1 vccd1 vccd1 op_cnt\[5\] sky130_fd_sc_hd__dfxtp_1
X_2865_ _0668_ u_bits.i_op1\[0\] _0675_ _0679_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__a31o_1
X_4604_ u_muldiv.o_div\[0\] u_muldiv.o_div\[1\] vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__nand2_1
X_5584_ clknet_leaf_38_i_clk _0231_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[1\] sky130_fd_sc_hd__dfxtp_1
X_4535_ _1999_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__clkbuf_1
X_2796_ _0490_ _0491_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__or2_1
X_4466_ u_muldiv.divisor\[59\] _1836_ _1946_ u_muldiv.divisor\[60\] _1961_ vssd1 vssd1
+ vccd1 vccd1 _0225_ sky130_fd_sc_hd__a221o_1
X_4397_ _1487_ u_bits.i_op2\[14\] _1899_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__or3_1
X_3417_ o_add[31] _1185_ _1186_ _1187_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__or4_4
X_3348_ _1133_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__nand2_4
X_3279_ _1015_ _1016_ _1074_ _1047_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__a211o_1
X_5018_ _2054_ _2370_ _2288_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_2650_ _0464_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__buf_2
X_4320_ _1842_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__buf_2
X_4251_ _1799_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
X_3202_ _0872_ _1002_ _0875_ _0871_ _0879_ _0923_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__mux4_1
X_4182_ u_wr_mux.i_reg_data2\[9\] i_reg_data2[9] _1756_ vssd1 vssd1 vccd1 vccd1 _1764_
+ sky130_fd_sc_hd__mux2_1
X_3133_ u_muldiv.dividend\[25\] _0742_ _0743_ u_muldiv.o_div\[25\] _0744_ vssd1 vssd1
+ vccd1 vccd1 _0938_ sky130_fd_sc_hd__a221o_1
X_3064_ _0871_ _0872_ _0696_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__mux2_1
X_3966_ i_rd[0] _1632_ _1636_ o_rd[0] vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__a22o_1
X_5705_ clknet_leaf_30_i_clk _0348_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_2917_ _0731_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__buf_2
X_3897_ _1255_ i_op1[2] _1599_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__mux2_1
X_5636_ clknet_leaf_42_i_clk _0283_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_2848_ _0533_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__clkbuf_4
X_2779_ _0592_ _0593_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__xnor2_4
X_5567_ clknet_leaf_8_i_clk _0214_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_4518_ u_muldiv.mul\[18\] u_muldiv.mul\[19\] _1989_ vssd1 vssd1 vccd1 vccd1 _1991_
+ sky130_fd_sc_hd__mux2_1
X_5498_ clknet_leaf_43_i_clk _0146_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_4449_ u_bits.i_op2\[25\] _1947_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__nand2_1
X_3820_ u_muldiv.dividend\[17\] _0721_ _0723_ u_muldiv.o_div\[17\] _0724_ vssd1 vssd1
+ vccd1 vccd1 _1540_ sky130_fd_sc_hd__a221o_1
X_3751_ _1110_ _1033_ _1473_ _1248_ _1475_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__a221o_1
X_2702_ _0457_ _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__xnor2_1
X_3682_ _1274_ _1410_ _1411_ _0624_ _1141_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__o32a_1
X_2633_ u_mux.i_group_mux vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__buf_2
X_5421_ clknet_leaf_52_i_clk _0069_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[12\] sky130_fd_sc_hd__dfxtp_4
X_5352_ _2009_ _2628_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__nor2_1
X_4303_ u_muldiv.i_on_end vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__clkinv_2
X_5283_ _2164_ _2606_ _2612_ _2613_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__a31o_1
X_4234_ csr_data\[0\] i_csr_data[0] _1789_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__mux2_1
X_4165_ o_wdata[1] i_reg_data2[1] _1745_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__mux2_1
X_3116_ _0825_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__clkbuf_4
X_4096_ _1720_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__clkbuf_1
X_3047_ u_muldiv.dividend\[23\] _0633_ _0722_ u_muldiv.o_div\[23\] _0724_ vssd1 vssd1
+ vccd1 vccd1 _0856_ sky130_fd_sc_hd__a221o_1
X_4998_ _1208_ _2345_ _2346_ _2353_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__a31o_1
X_3949_ _0996_ i_op1[27] _1621_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__mux2_1
X_5619_ clknet_leaf_45_i_clk _0266_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_16_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4921_ u_muldiv.quotient_msk\[28\] _2284_ _2283_ u_muldiv.quotient_msk\[29\] vssd1
+ vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__a22o_1
X_4852_ _2208_ _2249_ _2250_ _2251_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__a31o_1
X_3803_ _1333_ csr_data\[15\] _0731_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__o21ai_1
X_4783_ _1880_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__clkbuf_4
X_3734_ u_bits.i_op2\[11\] _1251_ _0926_ _1459_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__o22a_1
X_3665_ u_bits.i_op2\[6\] _0786_ _1272_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__a21oi_1
X_5404_ clknet_leaf_51_i_clk _0052_ vssd1 vssd1 vccd1 vccd1 o_rd[2] sky130_fd_sc_hd__dfxtp_2
X_3596_ _0453_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__buf_2
X_5335_ _1128_ _1585_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__nor2_1
X_5266_ _2030_ _2131_ _2132_ _2133_ vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__a31o_1
X_4217_ _1782_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__clkbuf_1
X_5197_ _2535_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__clkbuf_1
X_4148_ _1746_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__clkbuf_1
X_4079_ _1594_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__buf_6
X_3450_ _1215_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__clkbuf_1
X_3381_ _1159_ _1160_ _0507_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__a21bo_1
X_5120_ _2458_ _2089_ _2087_ vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__o21a_1
X_5051_ _2402_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__clkbuf_1
X_4002_ u_bits.i_op2\[9\] _1406_ _1657_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__mux2_1
X_4904_ u_muldiv.quotient_msk\[14\] _2280_ _2281_ u_muldiv.quotient_msk\[15\] vssd1
+ vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__a22o_1
X_4835_ u_muldiv.quotient_msk\[21\] _2233_ _2229_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__mux2_1
X_4766_ u_muldiv.quotient_msk\[7\] _2179_ _2156_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__mux2_1
X_3717_ _1443_ _1315_ _0970_ _0824_ _0670_ _0643_ vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__mux4_1
X_4697_ u_muldiv.dividend\[23\] u_muldiv.divisor\[23\] vssd1 vssd1 vccd1 vccd1 _2120_
+ sky130_fd_sc_hd__and2b_1
X_3648_ _1249_ _1375_ _1379_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__a21oi_1
X_3579_ _0645_ _0646_ _0630_ _0768_ _0658_ _0659_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__mux4_1
X_5318_ u_muldiv.divisor\[30\] _1838_ _1843_ u_muldiv.divisor\[31\] vssd1 vssd1 vccd1
+ vccd1 _0421_ sky130_fd_sc_hd__a22o_1
X_5249_ _2582_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__clkbuf_1
X_2950_ _0657_ _0702_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__and2b_1
X_2881_ u_bits.i_op2\[2\] vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__buf_4
X_4620_ u_muldiv.dividend\[13\] u_muldiv.divisor\[13\] vssd1 vssd1 vccd1 vccd1 _2043_
+ sky130_fd_sc_hd__and2b_1
X_4551_ _1135_ _2006_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__nor2_1
X_4482_ u_muldiv.mul\[1\] u_muldiv.mul\[2\] _1584_ vssd1 vssd1 vccd1 vccd1 _1972_
+ sky130_fd_sc_hd__mux2_1
X_3502_ _1233_ o_add[0] vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__and2_1
X_3433_ u_muldiv.i_on_wait _1202_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__nand2_1
X_3364_ _0594_ _1143_ _0605_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__o21ai_2
X_5103_ u_bits.i_op1\[13\] u_bits.i_op1\[14\] _2428_ vssd1 vssd1 vccd1 vccd1 _2450_
+ sky130_fd_sc_hd__or3_2
X_3295_ _0628_ _1082_ _1089_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__or3_2
X_5034_ _1250_ _2385_ _2386_ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__and3_1
X_4818_ _2181_ _2222_ _2224_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__a21oi_1
X_5798_ clknet_leaf_39_i_clk _0440_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[46\] sky130_fd_sc_hd__dfxtp_1
X_4749_ _2164_ _2166_ _2169_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__a21oi_1
X_3080_ _0857_ _0888_ _0446_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__a21oi_2
X_3982_ _0909_ _1112_ _1639_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__mux2_1
X_5721_ clknet_leaf_25_i_clk _0364_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2933_ u_muldiv.mul\[21\] _0740_ _0741_ u_muldiv.mul\[53\] _0745_ vssd1 vssd1 vccd1
+ vccd1 _0746_ sky130_fd_sc_hd__a221o_1
X_5652_ clknet_leaf_10_i_clk _0296_ vssd1 vssd1 vccd1 vccd1 op_cnt\[4\] sky130_fd_sc_hd__dfxtp_1
X_2864_ u_bits.i_op2\[2\] _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__and2b_1
X_4603_ u_muldiv.o_div\[0\] u_muldiv.o_div\[1\] vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__or2_1
X_5583_ clknet_leaf_35_i_clk _0230_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[0\] sky130_fd_sc_hd__dfxtp_1
X_2795_ _0488_ _0609_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__nand2_1
X_4534_ u_muldiv.mul\[26\] u_muldiv.mul\[27\] _1989_ vssd1 vssd1 vccd1 vccd1 _1999_
+ sky130_fd_sc_hd__mux2_1
X_4465_ _1959_ _1960_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__nor2_1
X_3416_ o_add[29] o_add[30] vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__or2_1
X_4396_ u_muldiv.divisor\[45\] _1867_ _1887_ u_muldiv.divisor\[46\] _1905_ vssd1 vssd1
+ vccd1 vccd1 _0211_ sky130_fd_sc_hd__a221o_1
X_3347_ _1131_ _1132_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__or2_1
X_5017_ _2054_ _2370_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__or2_1
X_3278_ _1023_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__inv_2
X_4250_ csr_data\[8\] i_csr_data[8] _1789_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__mux2_1
X_4181_ _1763_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__clkbuf_1
X_3201_ _1001_ _0944_ _0774_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__mux2_1
X_3132_ _0936_ _0937_ vssd1 vssd1 vccd1 vccd1 o_add[25] sky130_fd_sc_hd__xnor2_4
X_3063_ _0773_ _0781_ _0533_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__mux2_1
X_3965_ i_reg_write _1632_ _1636_ o_reg_write vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__a22o_1
X_5704_ clknet_leaf_30_i_clk _0347_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_2916_ _0730_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__inv_2
X_3896_ _1595_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__clkbuf_4
X_2847_ u_bits.i_op1\[10\] u_bits.i_op1\[9\] _0649_ vssd1 vssd1 vccd1 vccd1 _0662_
+ sky130_fd_sc_hd__mux2_1
X_5635_ clknet_leaf_41_i_clk _0282_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_2778_ u_bits.i_op1\[9\] u_muldiv.add_prev\[9\] _0450_ vssd1 vssd1 vccd1 vccd1 _0593_
+ sky130_fd_sc_hd__mux2_2
X_5566_ clknet_leaf_8_i_clk _0213_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_4517_ _1990_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__clkbuf_1
X_5497_ clknet_leaf_43_i_clk _0145_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_4448_ _0905_ _1942_ _1846_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__o21ai_1
X_4379_ _1445_ _1888_ _1846_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__o21a_1
X_3750_ u_bits.i_op2\[12\] _0777_ _0926_ _1474_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__o22a_1
X_2701_ _0460_ u_bits.i_op2\[12\] u_bits.i_op1\[12\] _0464_ vssd1 vssd1 vccd1 vccd1
+ _0516_ sky130_fd_sc_hd__a22o_1
X_3681_ _1406_ _1258_ _1272_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__a21oi_1
X_2632_ _0446_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__clkbuf_4
X_5420_ clknet_leaf_52_i_clk _0068_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[11\] sky130_fd_sc_hd__dfxtp_4
X_5351_ _1176_ _2628_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__nor2_1
X_4302_ u_muldiv.on_wait vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__clkbuf_4
X_5282_ u_muldiv.dividend\[31\] _2157_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__and2_1
X_4233_ i_to_trap _1638_ _1635_ o_to_trap vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__a22o_1
X_4164_ _1754_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__clkbuf_1
X_4095_ u_pc_sel.i_pc_next\[8\] i_pc_next[8] _1712_ vssd1 vssd1 vccd1 vccd1 _1720_
+ sky130_fd_sc_hd__mux2_1
X_3115_ _0904_ _0692_ _0691_ _0768_ _0658_ _0659_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__mux4_1
X_3046_ _0855_ vssd1 vssd1 vccd1 vccd1 o_add[23] sky130_fd_sc_hd__inv_2
X_4997_ _1207_ _2352_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__nor2_1
X_3948_ _1626_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__clkbuf_1
X_3879_ o_add[29] _1579_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__and2_1
X_5618_ clknet_leaf_45_i_clk _0265_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_5549_ clknet_leaf_6_i_clk mul_op2_signed_next vssd1 vssd1 vccd1 vccd1 u_muldiv.i_op2_signed
+ sky130_fd_sc_hd__dfxtp_1
X_4920_ u_muldiv.quotient_msk\[27\] _2284_ _2283_ u_muldiv.quotient_msk\[28\] vssd1
+ vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__a22o_1
X_4851_ u_muldiv.quotient_msk\[24\] u_muldiv.o_div\[24\] _1840_ vssd1 vssd1 vccd1
+ vccd1 _2251_ sky130_fd_sc_hd__o21a_1
X_3802_ _1331_ _1520_ _1522_ _1523_ _0728_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__o221a_1
X_4782_ u_muldiv.o_div\[10\] _2171_ _2195_ _2164_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__a22o_1
X_3733_ u_bits.i_op2\[11\] _1251_ _1267_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__a21oi_1
X_3664_ _1249_ _1391_ _1394_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__a21oi_1
X_5403_ clknet_leaf_51_i_clk _0051_ vssd1 vssd1 vccd1 vccd1 o_rd[1] sky130_fd_sc_hd__dfxtp_2
X_3595_ _0748_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__buf_2
X_5334_ _1130_ _1585_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__nor2_1
X_5265_ _2375_ _2135_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__nor2_1
X_5196_ u_muldiv.dividend\[23\] _2534_ _2485_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__mux2_1
X_4216_ u_wr_mux.i_reg_data2\[25\] i_reg_data2[25] _1778_ vssd1 vssd1 vccd1 vccd1
+ _1782_ sky130_fd_sc_hd__mux2_1
X_4147_ _0620_ i_funct3[0] _1745_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__mux2_1
X_4078_ u_bits.i_op2\[30\] _1639_ _1635_ _1710_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__a31o_1
X_3029_ _0677_ _0839_ _0779_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__mux2_1
X_3380_ _0577_ _1153_ _0521_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__o21ai_2
X_5050_ u_muldiv.dividend\[10\] _2401_ _2378_ vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__mux2_1
X_4001_ _1198_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__clkbuf_4
X_4903_ u_muldiv.quotient_msk\[13\] _2280_ _2281_ u_muldiv.quotient_msk\[14\] vssd1
+ vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__a22o_1
X_4834_ u_muldiv.o_div\[21\] _2170_ _2233_ _2196_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__a31o_1
X_4765_ _2165_ u_muldiv.o_div\[7\] _2179_ _1913_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__a31o_1
X_3716_ _1306_ _1309_ _0760_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__mux2_1
X_4696_ _2112_ _2118_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_15_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3647_ _1265_ _0797_ _1378_ _0634_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__o211ai_1
X_3578_ _1306_ _1309_ _1311_ _1312_ _0789_ _0674_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__mux4_1
X_5317_ u_muldiv.divisor\[29\] _1838_ _1843_ u_muldiv.divisor\[30\] vssd1 vssd1 vccd1
+ vccd1 _0420_ sky130_fd_sc_hd__a22o_1
X_5248_ u_muldiv.dividend\[28\] _2581_ _2485_ vssd1 vssd1 vccd1 vccd1 _2582_ sky130_fd_sc_hd__mux2_1
X_5179_ _0768_ _2511_ _2385_ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__o21ai_1
X_2880_ _0669_ _0690_ _0694_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__a21oi_1
X_4550_ _1137_ _2006_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__nor2_1
X_4481_ _1971_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__clkbuf_1
X_3501_ _0619_ o_add[1] vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__and2b_1
X_3432_ _1199_ _1201_ op_cnt\[0\] vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__a21oi_1
X_3363_ _1147_ vssd1 vssd1 vccd1 vccd1 o_add[8] sky130_fd_sc_hd__inv_2
X_5102_ _2447_ _2448_ vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__xnor2_1
X_3294_ _0925_ _1084_ _1085_ _0914_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__a221o_1
X_5033_ u_bits.i_op1\[7\] u_bits.i_op1\[8\] _2363_ vssd1 vssd1 vccd1 vccd1 _2386_
+ sky130_fd_sc_hd__or3_2
X_4817_ _2161_ _2223_ u_muldiv.o_div\[17\] vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__a21oi_1
X_5797_ clknet_leaf_39_i_clk _0439_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[45\] sky130_fd_sc_hd__dfxtp_1
X_4748_ _2167_ _2168_ u_muldiv.o_div\[3\] vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__a21oi_1
X_4679_ _2036_ _2038_ _2098_ _2101_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__a31o_1
X_3981_ _1641_ _1642_ _1643_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__a21o_1
X_2932_ u_muldiv.dividend\[21\] _0742_ _0743_ u_muldiv.o_div\[21\] _0744_ vssd1 vssd1
+ vccd1 vccd1 _0745_ sky130_fd_sc_hd__a221o_1
X_5720_ clknet_leaf_25_i_clk _0363_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_5651_ clknet_leaf_10_i_clk _0295_ vssd1 vssd1 vccd1 vccd1 op_cnt\[3\] sky130_fd_sc_hd__dfxtp_1
X_2863_ _0676_ _0677_ _0533_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__mux2_1
X_4602_ op_cnt\[5\] _2023_ _2025_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__o21a_1
X_5582_ clknet_leaf_36_i_clk _0229_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_2794_ _0493_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__inv_2
X_4533_ _1998_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__clkbuf_1
X_4464_ u_bits.i_op2\[28\] _1852_ _1958_ _1856_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__a31o_1
X_3415_ _0993_ _1024_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__nand2_1
X_4395_ _1832_ _1904_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__nor2_1
X_3346_ _1135_ vssd1 vssd1 vccd1 vccd1 o_add[5] sky130_fd_sc_hd__inv_2
X_5016_ _2055_ _2075_ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__or2_1
X_3277_ _1045_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__inv_2
X_4180_ u_wr_mux.i_reg_data2\[8\] i_reg_data2[8] _1756_ vssd1 vssd1 vccd1 vccd1 _1763_
+ sky130_fd_sc_hd__mux2_1
X_3200_ u_bits.i_op1\[27\] _0689_ _0778_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__mux2_1
X_3131_ _0898_ _0899_ _0901_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__a21bo_1
X_3062_ _0870_ _0772_ _0533_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__mux2_1
X_3964_ i_store _1632_ _1636_ o_store vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__a22o_1
X_5703_ clknet_leaf_30_i_clk _0346_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_2915_ o_res_src[1] vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__buf_2
X_3895_ _1598_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__clkbuf_1
X_2846_ u_bits.i_op1\[12\] u_bits.i_op1\[11\] _0657_ vssd1 vssd1 vccd1 vccd1 _0661_
+ sky130_fd_sc_hd__mux2_1
X_5634_ clknet_leaf_41_i_clk _0281_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_2777_ _0457_ _0591_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__xnor2_4
X_5565_ clknet_leaf_8_i_clk _0212_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_4516_ u_muldiv.mul\[17\] u_muldiv.mul\[18\] _1989_ vssd1 vssd1 vccd1 vccd1 _1990_
+ sky130_fd_sc_hd__mux2_1
X_5496_ clknet_leaf_43_i_clk _0144_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_4447_ _1841_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__buf_4
X_4378_ u_muldiv.divisor\[41\] _1867_ _1887_ u_muldiv.divisor\[42\] _1891_ vssd1 vssd1
+ vccd1 vccd1 _0207_ sky130_fd_sc_hd__a221o_1
X_3329_ _0749_ o_add[31] _1120_ _1121_ _0453_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__a221o_1
X_2700_ _0513_ _0514_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__nor2_1
X_3680_ _1249_ _1405_ _1409_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__a21oi_1
X_2631_ csr_read vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__buf_4
X_5350_ _2629_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__clkbuf_1
X_5281_ _2303_ _2609_ _2611_ _2165_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__a211o_1
X_4301_ i_inst_branch i_funct3[0] _1632_ _1825_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__a31o_1
X_4232_ _1790_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_1
X_4163_ o_wdata[0] i_reg_data2[0] _1745_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__mux2_1
X_3114_ _0916_ _0918_ _0919_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__a2bb2o_1
X_4094_ _1719_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__clkbuf_1
X_3045_ _0853_ _0854_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__xnor2_2
X_4996_ _2347_ _2349_ _2351_ _1826_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__o22a_1
X_3947_ _0689_ i_op1[26] _1621_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__mux2_1
X_3878_ _1024_ _1585_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__nor2_1
X_5617_ clknet_leaf_45_i_clk _0264_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2829_ _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__clkbuf_4
X_5548_ clknet_leaf_5_i_clk _0196_ vssd1 vssd1 vccd1 vccd1 u_adder.i_cmp_inverse sky130_fd_sc_hd__dfxtp_1
X_5479_ clknet_leaf_6_i_clk _0127_ vssd1 vssd1 vccd1 vccd1 alu_ctrl\[2\] sky130_fd_sc_hd__dfxtp_1
X_4850_ u_muldiv.o_div\[23\] u_muldiv.o_div\[24\] _2241_ vssd1 vssd1 vccd1 vccd1 _2250_
+ sky130_fd_sc_hd__or3_2
X_3801_ u_muldiv.mul\[15\] _0748_ _1400_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__o21ai_1
X_4781_ _2165_ _2193_ _2194_ _1842_ u_muldiv.quotient_msk\[10\] vssd1 vssd1 vccd1
+ vccd1 _2195_ sky130_fd_sc_hd__a32o_1
X_3732_ _1457_ _1344_ _0998_ _0824_ _0707_ _0643_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__mux4_1
X_3663_ _0674_ _1110_ _0841_ _1393_ _0858_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__a311o_1
X_5402_ clknet_leaf_51_i_clk _0050_ vssd1 vssd1 vccd1 vccd1 o_rd[0] sky130_fd_sc_hd__dfxtp_2
X_3594_ u_muldiv.mul\[34\] _1325_ _1328_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__a21oi_1
X_5333_ _2627_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__clkbuf_1
X_5264_ _0699_ _2362_ _2594_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__nand3_1
X_5195_ _1208_ _2525_ _2526_ _2533_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__a31o_1
X_4215_ _1781_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__clkbuf_1
X_4146_ _1711_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__buf_6
X_4077_ u_bits.i_op2\[31\] _1634_ _1596_ i_op2[31] vssd1 vssd1 vccd1 vccd1 _1710_
+ sky130_fd_sc_hd__a22o_1
X_3028_ _0658_ u_bits.i_op1\[0\] vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__and2b_1
X_4979_ u_muldiv.dividend\[5\] u_muldiv.dividend\[4\] _2315_ vssd1 vssd1 vccd1 vccd1
+ _2336_ sky130_fd_sc_hd__or3_1
X_4000_ _1641_ _1655_ _1656_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__a21o_1
X_4902_ u_muldiv.quotient_msk\[12\] _2280_ _2281_ u_muldiv.quotient_msk\[13\] vssd1
+ vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__a22o_1
X_4833_ _2236_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__clkbuf_1
X_4764_ _2154_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__buf_2
X_3715_ _1441_ _1442_ _1336_ u_pc_sel.i_pc_next\[9\] vssd1 vssd1 vccd1 vccd1 o_result[9]
+ sky130_fd_sc_hd__a2bb2o_2
X_4695_ _2113_ _2117_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__nand2_1
X_3646_ _1376_ _1257_ _1293_ _1377_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__a2bb2o_1
X_3577_ _0786_ _1258_ _0785_ _1250_ _0651_ _0774_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__mux4_1
X_5316_ u_muldiv.divisor\[28\] _1838_ _2617_ u_muldiv.divisor\[29\] vssd1 vssd1 vccd1
+ vccd1 _0419_ sky130_fd_sc_hd__a22o_1
X_5247_ _2575_ _2579_ _1877_ _2580_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__o2bb2a_1
X_5178_ _2104_ _2035_ _2102_ _1839_ vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__a31o_1
X_4129_ _1736_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__clkbuf_1
X_3500_ _1192_ u_wr_mux.i_reg_data2\[31\] _1241_ vssd1 vssd1 vccd1 vccd1 o_wdata[31]
+ sky130_fd_sc_hd__a21o_2
X_4480_ u_muldiv.mul\[0\] u_muldiv.mul\[1\] _1584_ vssd1 vssd1 vccd1 vccd1 _1971_
+ sky130_fd_sc_hd__mux2_1
X_3431_ _1198_ op_cnt\[5\] _1200_ op_cnt\[4\] vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__or4b_1
X_3362_ _1143_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__nand2_2
X_5101_ _2039_ _2082_ vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__and2b_1
X_3293_ _0699_ u_bits.i_op2\[30\] _0636_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__o22a_1
X_5032_ _2292_ vssd1 vssd1 vccd1 vccd1 _2385_ sky130_fd_sc_hd__buf_2
X_4816_ u_muldiv.quotient_msk\[17\] _2218_ _2156_ vssd1 vssd1 vccd1 vccd1 _2223_ sky130_fd_sc_hd__mux2_1
X_5796_ clknet_leaf_34_i_clk _0438_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[44\] sky130_fd_sc_hd__dfxtp_1
X_4747_ u_muldiv.quotient_msk\[3\] _2158_ _2156_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__mux2_1
X_4678_ _2034_ _2100_ _2032_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__or3b_1
X_3629_ _0751_ _0708_ _1361_ _0710_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_14_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3980_ _1112_ _1637_ _1638_ i_op2[1] vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__a22o_1
X_2931_ _0724_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__clkbuf_4
X_5650_ clknet_leaf_11_i_clk _0294_ vssd1 vssd1 vccd1 vccd1 op_cnt\[2\] sky130_fd_sc_hd__dfxtp_1
X_4601_ op_cnt\[5\] _2023_ _1204_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__a21oi_1
X_2862_ u_bits.i_op1\[2\] u_bits.i_op1\[1\] _0656_ vssd1 vssd1 vccd1 vccd1 _0677_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_29_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2793_ _0579_ _0607_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__or2_1
X_5581_ clknet_leaf_3_i_clk _0228_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_4532_ u_muldiv.mul\[25\] u_muldiv.mul\[26\] _1989_ vssd1 vssd1 vccd1 vccd1 _1998_
+ sky130_fd_sc_hd__mux2_1
X_4463_ _1868_ _1958_ u_bits.i_op2\[28\] vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__a21oi_1
X_3414_ o_add[25] o_add[26] _1183_ _1184_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__or4_1
X_4394_ u_bits.i_op2\[14\] _1903_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__xnor2_1
X_3345_ _0566_ _1134_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__xor2_4
X_3276_ _1070_ _1071_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__nand2_2
X_5015_ u_muldiv.dividend\[8\] _2361_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__xor2_1
X_5779_ clknet_leaf_21_i_clk _0422_ vssd1 vssd1 vccd1 vccd1 u_muldiv.outsign sky130_fd_sc_hd__dfxtp_2
X_3130_ _0934_ _0935_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__xnor2_4
X_3061_ u_bits.i_op1\[23\] u_bits.i_op1\[22\] _0649_ vssd1 vssd1 vccd1 vccd1 _0870_
+ sky130_fd_sc_hd__mux2_1
X_3963_ _1635_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__buf_2
X_5702_ clknet_leaf_30_i_clk _0345_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_2914_ _0728_ csr_data\[20\] vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__or2_1
X_3894_ _0791_ i_op1[1] _1596_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__mux2_1
X_5633_ clknet_leaf_42_i_clk _0280_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_2845_ _0653_ _0654_ _0655_ u_bits.i_op1\[13\] _0658_ _0659_ vssd1 vssd1 vccd1 vccd1
+ _0660_ sky130_fd_sc_hd__mux4_1
X_5564_ clknet_leaf_3_i_clk _0211_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_4515_ _1583_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__clkbuf_4
X_2776_ _0460_ u_bits.i_op2\[9\] u_bits.i_op1\[9\] _0464_ vssd1 vssd1 vccd1 vccd1
+ _0591_ sky130_fd_sc_hd__a22o_1
X_5495_ clknet_leaf_43_i_clk _0143_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_4446_ u_muldiv.divisor\[55\] _1878_ _1829_ u_muldiv.divisor\[56\] _1945_ vssd1 vssd1
+ vccd1 vccd1 _0221_ sky130_fd_sc_hd__o221a_1
X_4377_ _1889_ _1890_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__nor2_1
X_3328_ _0629_ _1115_ _0955_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__a21oi_1
X_3259_ _0697_ u_bits.i_op1\[28\] _0778_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__mux2_1
X_5280_ _0620_ _2610_ _2375_ _0702_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__o211a_1
X_4300_ _1171_ _1638_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__nor2_1
X_4231_ _0446_ i_csr_read _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__mux2_1
X_4162_ _1753_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__clkbuf_1
X_3113_ _0673_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__buf_4
X_4093_ u_pc_sel.i_pc_next\[7\] i_pc_next[7] _1712_ vssd1 vssd1 vccd1 vccd1 _1719_
+ sky130_fd_sc_hd__mux2_1
X_3044_ _0812_ _0815_ _0810_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__a21bo_1
X_4995_ _0786_ _2350_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__xnor2_1
X_3946_ _1625_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__clkbuf_1
X_3877_ _0993_ _1585_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__nor2_1
X_5616_ clknet_leaf_44_i_clk _0263_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2828_ _0642_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__clkbuf_4
X_5547_ clknet_leaf_11_i_clk _0195_ vssd1 vssd1 vccd1 vccd1 csr_data\[31\] sky130_fd_sc_hd__dfxtp_1
X_2759_ _0571_ _0572_ _0573_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__o21a_1
X_5478_ clknet_leaf_46_i_clk _0126_ vssd1 vssd1 vccd1 vccd1 u_mux.i_group_mux sky130_fd_sc_hd__dfxtp_2
X_4429_ u_bits.i_op2\[21\] _1931_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__xnor2_1
X_4780_ u_muldiv.o_div\[9\] u_muldiv.o_div\[10\] _2186_ vssd1 vssd1 vccd1 vccd1 _2194_
+ sky130_fd_sc_hd__or3_1
X_3800_ u_muldiv.mul\[47\] _0741_ _1521_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__a21oi_1
X_3731_ _1337_ _1339_ _0760_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__mux2_1
X_3662_ u_bits.i_op2\[6\] _0786_ _0926_ _1392_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__o22a_1
X_3593_ u_muldiv.dividend\[2\] _1326_ _1327_ u_muldiv.o_div\[2\] _0717_ vssd1 vssd1
+ vccd1 vccd1 _1328_ sky130_fd_sc_hd__a221o_1
X_5401_ clknet_leaf_51_i_clk _0049_ vssd1 vssd1 vccd1 vccd1 o_reg_write sky130_fd_sc_hd__dfxtp_2
X_5332_ o_add[1] _1579_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__and2_1
X_5263_ _2362_ _2594_ _0699_ vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__a21o_1
X_5194_ _2375_ _2527_ _2529_ _2532_ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__o31a_1
X_4214_ u_wr_mux.i_reg_data2\[24\] i_reg_data2[24] _1778_ vssd1 vssd1 vccd1 vccd1
+ _1781_ sky130_fd_sc_hd__mux2_1
X_4145_ _1744_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__clkbuf_1
X_4076_ _1689_ _1708_ _1709_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__a21o_1
X_3027_ _0666_ _0676_ _0659_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__mux2_1
X_4978_ u_muldiv.dividend\[4\] _2315_ u_muldiv.dividend\[5\] vssd1 vssd1 vccd1 vccd1
+ _2335_ sky130_fd_sc_hd__o21ai_1
X_3929_ _1616_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__clkbuf_1
X_4901_ u_muldiv.quotient_msk\[11\] _2280_ _2281_ u_muldiv.quotient_msk\[12\] vssd1
+ vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__a22o_1
X_4832_ u_muldiv.o_div\[20\] _2235_ _2154_ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__mux2_1
X_4763_ u_muldiv.o_div\[6\] _2171_ _2180_ _2164_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__a22o_1
X_4694_ _2116_ vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__inv_2
X_3714_ _1333_ csr_data\[9\] _1388_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__o21ai_1
X_3645_ _1376_ _1257_ _0867_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__a21o_1
X_3576_ _1255_ _0794_ _1310_ _1257_ _0651_ _1112_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__mux4_1
X_5315_ u_muldiv.divisor\[27\] _1838_ _2617_ u_muldiv.divisor\[28\] vssd1 vssd1 vccd1
+ vccd1 _0418_ sky130_fd_sc_hd__a22o_1
X_5246_ u_muldiv.dividend\[28\] _2564_ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__xor2_1
X_5177_ _2517_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__clkbuf_1
X_4128_ o_pc_target[7] i_pc_target[7] _1734_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__mux2_1
X_4059_ u_bits.i_op2\[26\] _0905_ _1681_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__mux2_1
X_3430_ op_cnt\[1\] op_cnt\[2\] op_cnt\[3\] vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__nand3_1
X_3361_ _0568_ _0576_ _0598_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__nand3_1
X_5100_ _2040_ _2436_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__nand2_1
X_5031_ _2382_ _2383_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__xnor2_1
X_3292_ _0617_ _0638_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__and3_1
X_4815_ _2170_ u_muldiv.o_div\[17\] _2218_ _2196_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__a31o_1
X_5795_ clknet_leaf_37_i_clk _0437_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[43\] sky130_fd_sc_hd__dfxtp_1
X_4746_ _2153_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__clkbuf_4
X_4677_ _2033_ _2099_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__nand2_1
X_3628_ _0687_ _1360_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__nor2_1
X_3559_ _1112_ _0791_ _1293_ _1294_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__a2bb2o_1
X_5229_ u_muldiv.dividend\[27\] u_muldiv.dividend\[26\] _2552_ vssd1 vssd1 vccd1 vccd1
+ _2564_ sky130_fd_sc_hd__or3_1
X_2930_ _0722_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__buf_2
X_4600_ op_cnt\[4\] _2021_ _2024_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__o21a_1
X_2861_ u_bits.i_op1\[4\] u_bits.i_op1\[3\] _0656_ vssd1 vssd1 vccd1 vccd1 _0676_
+ sky130_fd_sc_hd__mux2_1
X_5580_ clknet_leaf_9_i_clk _0227_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_2792_ _0602_ _0603_ _0590_ _0605_ _0606_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__o221a_1
X_4531_ _1997_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkbuf_1
X_4462_ u_bits.i_op2\[26\] u_bits.i_op2\[27\] _1942_ _1951_ vssd1 vssd1 vccd1 vccd1
+ _1958_ sky130_fd_sc_hd__or4_1
X_3413_ _0855_ _0903_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__nand2_1
X_4393_ _1487_ _1899_ _1845_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__o21a_1
X_3344_ _0571_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__nand2_1
X_3275_ _1068_ _1069_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__or2_1
X_5014_ _2157_ _2359_ _2367_ _2368_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__o31a_1
X_5778_ clknet_leaf_8_i_clk _0421_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_4729_ _1839_ _2135_ _2138_ _2151_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__o31a_4
X_3060_ _0692_ u_bits.i_op2\[23\] _0636_ _0868_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__o22a_1
X_5701_ clknet_leaf_29_i_clk _0344_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_3962_ _1204_ _1634_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__nor2_4
X_2913_ csr_read vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__clkinv_4
X_3893_ _1597_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__clkbuf_1
X_5632_ clknet_leaf_42_i_clk _0279_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_2844_ _0533_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__clkbuf_4
X_5563_ clknet_leaf_5_i_clk _0210_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_4514_ _1988_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__clkbuf_1
X_2775_ _0584_ _0589_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__nand2_1
X_5494_ clknet_leaf_43_i_clk _0142_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4445_ _0905_ _1943_ _1944_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__o21ai_1
X_4376_ _1445_ _1852_ _1888_ _1856_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__a31o_1
X_3327_ _0914_ _1109_ _1119_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__a21o_1
X_3258_ _0920_ _1053_ _1054_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__a21bo_1
X_3189_ _0989_ _0990_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_13_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_28_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4230_ _1711_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__clkbuf_4
X_4161_ _1274_ i_alu_ctrl[4] _1745_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__mux2_1
X_4092_ _1718_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__clkbuf_1
X_3112_ _0667_ _0678_ _0758_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__mux2_1
X_3043_ _0851_ _0852_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__nor2_1
X_4994_ _1310_ _1257_ _2328_ _2292_ vssd1 vssd1 vccd1 vccd1 _2350_ sky130_fd_sc_hd__o31a_1
X_3945_ _0943_ i_op1[25] _1621_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__mux2_1
X_5615_ clknet_leaf_46_i_clk _0262_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3876_ _1587_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__clkbuf_1
X_2827_ u_bits.i_op2\[4\] vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__clkbuf_4
X_5546_ clknet_leaf_11_i_clk _0194_ vssd1 vssd1 vccd1 vccd1 csr_data\[30\] sky130_fd_sc_hd__dfxtp_1
X_2758_ _0564_ _0565_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__nand2_1
X_5477_ clknet_leaf_48_i_clk _0125_ vssd1 vssd1 vccd1 vccd1 u_muldiv.i_is_div sky130_fd_sc_hd__dfxtp_1
X_2689_ _0448_ u_bits.i_op1\[14\] _0497_ _0503_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__a31o_1
X_4428_ u_bits.i_op2\[20\] _1927_ _1845_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__o21a_1
X_4359_ _1874_ _1875_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__nor2_1
X_3730_ _1455_ _1456_ _1336_ u_pc_sel.i_pc_next\[10\] vssd1 vssd1 vccd1 vccd1 o_result[10]
+ sky130_fd_sc_hd__a2bb2o_2
X_3661_ u_bits.i_op2\[6\] _0786_ _0867_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__a21oi_1
X_3592_ _0722_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__buf_2
X_5400_ clknet_leaf_1_i_clk _0048_ vssd1 vssd1 vccd1 vccd1 o_store sky130_fd_sc_hd__dfxtp_2
X_5331_ _2626_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__clkbuf_1
X_5262_ _0996_ _1029_ _0697_ _2568_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__or4_1
X_5193_ _2288_ _2531_ _1206_ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__a21oi_1
X_4213_ _1780_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__clkbuf_1
X_4144_ o_pc_target[15] i_pc_target[15] _1734_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__mux2_1
X_4075_ u_bits.i_op2\[30\] _1634_ _1596_ i_op2[30] vssd1 vssd1 vccd1 vccd1 _1709_
+ sky130_fd_sc_hd__a22o_1
X_3026_ _0832_ _0833_ _0835_ _0836_ _0825_ _0707_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__mux4_1
X_4977_ _2334_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__clkbuf_1
X_3928_ _0647_ i_op1[17] _1610_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__mux2_1
X_3859_ _0749_ o_add[19] _1575_ _1576_ _0453_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__a221o_1
X_5529_ clknet_leaf_15_i_clk _0177_ vssd1 vssd1 vccd1 vccd1 csr_data\[13\] sky130_fd_sc_hd__dfxtp_1
X_4900_ u_muldiv.quotient_msk\[10\] _2280_ _2281_ u_muldiv.quotient_msk\[11\] vssd1
+ vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__a22o_1
X_4831_ _2208_ _2232_ _2233_ _2234_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__a31o_1
X_4762_ _2165_ _2178_ _2179_ _1842_ u_muldiv.quotient_msk\[6\] vssd1 vssd1 vccd1 vccd1
+ _2180_ sky130_fd_sc_hd__a32o_1
X_4693_ _2114_ _2115_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__or2_1
X_3713_ _0454_ _1437_ _1439_ _1440_ _1357_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__o221a_1
X_3644_ u_bits.i_op2\[5\] vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_2_2__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3575_ u_bits.i_op1\[4\] vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__buf_4
X_5314_ u_muldiv.divisor\[26\] _1838_ _2617_ u_muldiv.divisor\[27\] vssd1 vssd1 vccd1
+ vccd1 _0417_ sky130_fd_sc_hd__a22o_1
X_5245_ _1827_ _2577_ _2578_ _1840_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__a31o_1
X_5176_ u_muldiv.dividend\[21\] _2516_ _2485_ vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__mux2_1
X_4127_ _1735_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__clkbuf_1
X_4058_ _1689_ _1696_ _1697_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__a21o_1
X_3009_ _0533_ _0819_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__and2b_1
X_3360_ _1145_ vssd1 vssd1 vccd1 vccd1 o_add[9] sky130_fd_sc_hd__inv_2
X_5030_ _2051_ _2076_ vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__and2b_1
X_3291_ _0699_ u_bits.i_op2\[30\] vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__nand2_2
X_4814_ _2221_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__clkbuf_1
X_5794_ clknet_leaf_35_i_clk _0436_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[42\] sky130_fd_sc_hd__dfxtp_1
X_4745_ _2165_ u_muldiv.o_div\[3\] _2158_ _1913_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__a31o_1
X_4676_ u_muldiv.dividend\[20\] u_muldiv.divisor\[20\] vssd1 vssd1 vccd1 vccd1 _2099_
+ sky130_fd_sc_hd__or2b_1
X_3627_ _1253_ _1261_ _1259_ _1252_ _0760_ _0879_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__mux4_1
X_3558_ _1112_ _0791_ _0866_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__a21o_1
X_3489_ o_wdata[2] _1233_ _0799_ u_wr_mux.i_reg_data2\[10\] vssd1 vssd1 vccd1 vccd1
+ _1236_ sky130_fd_sc_hd__a22o_1
X_5228_ _2563_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__clkbuf_1
X_5159_ _0646_ _2492_ _2385_ vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__o21ai_1
X_2860_ _0650_ _0663_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__nor2_1
X_2791_ _0582_ _0583_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__nand2_1
X_4530_ u_muldiv.mul\[24\] u_muldiv.mul\[25\] _1989_ vssd1 vssd1 vccd1 vccd1 _1997_
+ sky130_fd_sc_hd__mux2_1
X_4461_ u_muldiv.divisor\[58\] _1836_ _1946_ u_muldiv.divisor\[59\] _1957_ vssd1 vssd1
+ vccd1 vccd1 _0224_ sky130_fd_sc_hd__a221o_1
X_3412_ o_add[20] _1172_ _1173_ _1182_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__or4_1
X_4392_ u_muldiv.divisor\[44\] _1867_ _1887_ u_muldiv.divisor\[45\] _1902_ vssd1 vssd1
+ vccd1 vccd1 _0210_ sky130_fd_sc_hd__a221o_1
X_3343_ _1131_ _1132_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__nand2_2
X_3274_ _1068_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__nand2_4
X_5013_ u_muldiv.dividend\[7\] _2154_ vssd1 vssd1 vccd1 vccd1 _2368_ sky130_fd_sc_hd__or2_1
X_5777_ clknet_leaf_11_i_clk _0420_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_2989_ _0628_ _0767_ _0771_ _0801_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__or4_1
X_4728_ _1831_ _2150_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__nand2_1
X_4659_ u_muldiv.divisor\[15\] u_muldiv.dividend\[15\] vssd1 vssd1 vccd1 vccd1 _2082_
+ sky130_fd_sc_hd__or2b_1
X_3961_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__buf_2
X_5700_ clknet_leaf_29_i_clk _0343_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_2912_ _0454_ _0716_ _0726_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__o21a_1
X_3892_ _0917_ i_op1[0] _1596_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__mux2_1
X_2843_ _0657_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__buf_4
X_5631_ clknet_leaf_41_i_clk _0278_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_2774_ _0587_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__xor2_4
X_5562_ clknet_leaf_5_i_clk _0209_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_4513_ u_muldiv.mul\[16\] u_muldiv.mul\[17\] _1978_ vssd1 vssd1 vccd1 vccd1 _1988_
+ sky130_fd_sc_hd__mux2_1
X_5493_ clknet_leaf_50_i_clk _0141_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[11\]
+ sky130_fd_sc_hd__dfxtp_4
X_4444_ _0905_ _1943_ _1832_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__a21oi_1
X_4375_ _1868_ _1888_ _1445_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__a21oi_1
X_3326_ _1110_ _1114_ _1118_ _0858_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_9_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3257_ _0760_ _0793_ _0796_ _0673_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__a211o_1
X_3188_ _0987_ _0988_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__nor2_1
X_4160_ _1752_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__clkbuf_1
X_3111_ _0707_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__nand2_1
X_4091_ u_pc_sel.i_pc_next\[6\] i_pc_next[6] _1712_ vssd1 vssd1 vccd1 vccd1 _1718_
+ sky130_fd_sc_hd__mux2_1
X_3042_ _0849_ _0850_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__nor2_1
X_4993_ _1826_ _2348_ vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__nand2_1
X_3944_ _1624_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__clkbuf_1
X_3875_ o_add[26] _1579_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__and2_1
X_5614_ clknet_leaf_44_i_clk _0261_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2826_ _0630_ u_bits.i_op2\[20\] _0637_ _0640_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__o22ai_1
X_5545_ clknet_leaf_11_i_clk _0193_ vssd1 vssd1 vccd1 vccd1 csr_data\[29\] sky130_fd_sc_hd__dfxtp_1
X_2757_ _0564_ _0565_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__nor2_1
X_5476_ clknet_leaf_23_i_clk _0124_ vssd1 vssd1 vccd1 vccd1 o_funct3[2] sky130_fd_sc_hd__dfxtp_4
X_2688_ u_mux.i_group_mux u_bits.i_op2\[14\] vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__and2b_1
X_4427_ u_muldiv.divisor\[51\] _1878_ _1833_ _1929_ _1930_ vssd1 vssd1 vccd1 vccd1
+ _0217_ sky130_fd_sc_hd__o221a_1
X_4358_ _1406_ _1850_ _1873_ _1856_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__a31o_1
X_4289_ _1819_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
X_3309_ _1101_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__nand2_1
X_3660_ _1390_ _0826_ _0751_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__mux2_1
X_3591_ _0633_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__buf_2
X_5330_ o_add[0] _1579_ vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__and2_1
X_5261_ _2593_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__clkbuf_1
X_4212_ u_wr_mux.i_reg_data2\[23\] i_reg_data2[23] _1778_ vssd1 vssd1 vccd1 vccd1
+ _1780_ sky130_fd_sc_hd__mux2_1
X_5192_ _0692_ _2530_ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__xnor2_1
X_4143_ _1743_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__clkbuf_1
X_4074_ u_bits.i_op2\[31\] u_bits.i_op2\[29\] _1198_ vssd1 vssd1 vccd1 vccd1 _1708_
+ sky130_fd_sc_hd__mux2_1
X_3025_ _0662_ _0665_ _0779_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4976_ u_muldiv.dividend\[4\] _2333_ _2244_ vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__mux2_1
X_3927_ _1615_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__clkbuf_1
X_3858_ _0908_ _1569_ _0955_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_27_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3789_ _1510_ _1511_ _0730_ u_pc_sel.i_pc_next\[14\] vssd1 vssd1 vccd1 vccd1 o_result[14]
+ sky130_fd_sc_hd__a2bb2o_2
X_2809_ _0623_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__buf_2
X_5528_ clknet_leaf_13_i_clk _0176_ vssd1 vssd1 vccd1 vccd1 csr_data\[12\] sky130_fd_sc_hd__dfxtp_1
X_5459_ clknet_leaf_10_i_clk _0107_ vssd1 vssd1 vccd1 vccd1 o_pc_target[1] sky130_fd_sc_hd__dfxtp_2
X_4830_ u_muldiv.quotient_msk\[20\] u_muldiv.o_div\[20\] _1840_ vssd1 vssd1 vccd1
+ vccd1 _2234_ sky130_fd_sc_hd__o21a_1
X_4761_ u_muldiv.o_div\[5\] u_muldiv.o_div\[6\] _2173_ vssd1 vssd1 vccd1 vccd1 _2179_
+ sky130_fd_sc_hd__or3_1
X_4692_ u_muldiv.dividend\[26\] u_muldiv.divisor\[26\] vssd1 vssd1 vccd1 vccd1 _2115_
+ sky130_fd_sc_hd__and2b_1
X_3712_ u_muldiv.mul\[9\] _1330_ _1400_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__o21ai_1
X_3643_ _1374_ _0766_ _0751_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__mux2_1
X_5313_ u_muldiv.divisor\[25\] _2616_ _2617_ u_muldiv.divisor\[26\] vssd1 vssd1 vccd1
+ vccd1 _0416_ sky130_fd_sc_hd__a22o_1
X_3574_ _1307_ _1308_ _0779_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__mux2_1
X_5244_ _1029_ _2576_ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__or2_1
X_5175_ _1208_ _2506_ _2507_ _2515_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__a31o_1
X_4126_ o_pc_target[6] i_pc_target[6] _1734_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__mux2_1
X_4057_ _0905_ _1687_ _1675_ i_op2[24] vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__a22o_1
X_3008_ u_bits.i_op1\[26\] u_bits.i_op1\[27\] _0656_ vssd1 vssd1 vccd1 vccd1 _0819_
+ sky130_fd_sc_hd__mux2_1
X_4959_ _2059_ _2317_ vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__nand2_1
X_3290_ _0835_ _0836_ _0838_ _0840_ _0669_ _0670_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__mux4_1
X_4813_ u_muldiv.o_div\[16\] _2220_ _2154_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__mux2_1
X_5793_ clknet_leaf_35_i_clk _0435_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[41\] sky130_fd_sc_hd__dfxtp_1
X_4744_ _1208_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__clkbuf_4
X_4675_ _2039_ _2083_ _2095_ _2097_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__o31a_1
X_3626_ _1358_ _1359_ _1336_ u_pc_sel.i_pc_next\[3\] vssd1 vssd1 vccd1 vccd1 o_result[3]
+ sky130_fd_sc_hd__a2bb2o_2
X_3557_ _0620_ _0635_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__or2_1
X_5227_ u_muldiv.dividend\[26\] _2562_ _2485_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__mux2_1
X_3488_ _1192_ u_wr_mux.i_reg_data2\[25\] _1235_ vssd1 vssd1 vccd1 vccd1 o_wdata[25]
+ sky130_fd_sc_hd__a21o_2
X_5158_ _2499_ _2100_ vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__xor2_1
X_5089_ _2043_ _2081_ _2042_ vssd1 vssd1 vccd1 vccd1 _2437_ sky130_fd_sc_hd__o21a_1
X_4109_ _1727_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__clkbuf_1
X_2790_ _0592_ _0593_ _0604_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__o21ai_1
X_4460_ u_bits.i_op2\[27\] _1955_ _1956_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__o21a_1
X_3411_ o_add[12] o_add[16] _1177_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__or4b_1
X_4391_ _1900_ _1901_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__nor2_1
X_3342_ _0551_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__inv_2
X_3273_ u_bits.i_op1\[30\] u_muldiv.add_prev\[30\] _0452_ vssd1 vssd1 vccd1 vccd1
+ _1069_ sky130_fd_sc_hd__mux2_1
X_5012_ _1209_ _2360_ _2361_ _2366_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__a31o_1
X_5776_ clknet_leaf_11_i_clk _0419_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_2988_ _0672_ _0790_ _0798_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__o211a_1
X_4727_ _2146_ _2147_ _2148_ _2149_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__or4_1
X_4658_ _2046_ _2047_ _2079_ _2044_ _2080_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__o311a_1
X_3609_ _1287_ _0752_ _0659_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__mux2_1
X_4589_ _1204_ op_cnt\[0\] vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__nor2_1
X_3960_ i_flush i_reset_n vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__or2b_1
X_2911_ u_muldiv.mul\[20\] _0717_ _0720_ u_muldiv.mul\[52\] _0725_ vssd1 vssd1 vccd1
+ vccd1 _0726_ sky130_fd_sc_hd__a221o_1
X_3891_ _1595_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__clkbuf_4
X_2842_ _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__clkbuf_4
X_5630_ clknet_leaf_41_i_clk _0277_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_5561_ clknet_leaf_7_i_clk _0208_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_2773_ u_bits.i_op1\[10\] u_muldiv.add_prev\[10\] _0449_ vssd1 vssd1 vccd1 vccd1
+ _0588_ sky130_fd_sc_hd__mux2_2
X_4512_ _1987_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__clkbuf_1
X_5492_ clknet_leaf_50_i_clk _0140_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[10\]
+ sky130_fd_sc_hd__dfxtp_4
X_4443_ _1850_ _1942_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__nand2_1
X_4374_ u_bits.i_op2\[9\] _1883_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__or2_1
X_3325_ _0711_ _0860_ _0911_ _1117_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__a31o_1
X_3256_ _0780_ _0787_ _0758_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__mux2_1
X_3187_ _0987_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__and2_1
X_5759_ clknet_leaf_19_i_clk _0402_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_3110_ u_bits.i_op1\[0\] vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__buf_4
X_4090_ _1717_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__clkbuf_1
X_3041_ _0849_ _0850_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__and2_1
X_4992_ _2056_ _2071_ _2072_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__or3_1
X_3943_ _0904_ i_op1[24] _1621_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__mux2_1
X_3874_ _1586_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__clkbuf_1
X_5613_ clknet_leaf_34_i_clk _0260_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[30\] sky130_fd_sc_hd__dfxtp_1
X_2825_ _0618_ _0639_ _0631_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__and3_1
X_5544_ clknet_leaf_16_i_clk _0192_ vssd1 vssd1 vccd1 vccd1 csr_data\[28\] sky130_fd_sc_hd__dfxtp_1
X_2756_ _0549_ _0550_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__nand2_1
X_2687_ _0500_ _0501_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__nor2_1
X_5475_ clknet_leaf_6_i_clk _0123_ vssd1 vssd1 vccd1 vccd1 o_funct3[1] sky130_fd_sc_hd__dfxtp_4
X_4426_ u_muldiv.divisor\[52\] _1829_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__or2_1
X_4357_ _1868_ _1873_ _1406_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__a21oi_1
X_4288_ csr_data\[26\] i_csr_data[26] _1811_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__mux2_1
X_3308_ _1095_ _1100_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__or2_1
X_3239_ _1029_ u_bits.i_op2\[28\] _0634_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_8_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3590_ _0719_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__buf_2
X_5260_ u_muldiv.dividend\[29\] _2592_ _2485_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__mux2_1
X_4211_ _1779_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__clkbuf_1
X_5191_ _0768_ _0691_ _2511_ _2292_ vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__o31a_1
X_4142_ o_pc_target[14] i_pc_target[14] _1734_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__mux2_1
X_4073_ _1689_ _1706_ _1707_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__a21o_1
X_3024_ _0834_ _0661_ _0783_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__mux2_1
X_4975_ _2331_ _2332_ _2229_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__mux2_1
X_3926_ _0653_ i_op1[16] _1610_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__mux2_1
X_3857_ _0858_ _1568_ _1571_ _1574_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__or4_1
X_3788_ _1333_ csr_data\[14\] _1388_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__o21ai_1
X_2808_ u_mux.i_add_override _0622_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__nor2_2
X_5527_ clknet_leaf_13_i_clk _0175_ vssd1 vssd1 vccd1 vccd1 csr_data\[11\] sky130_fd_sc_hd__dfxtp_1
X_2739_ _0455_ _0553_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__xnor2_2
X_5458_ clknet_leaf_50_i_clk _0106_ vssd1 vssd1 vccd1 vccd1 o_res_src[2] sky130_fd_sc_hd__dfxtp_2
X_5389_ clknet_leaf_49_i_clk _0037_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[21\] sky130_fd_sc_hd__dfxtp_2
X_4409_ u_bits.i_op2\[17\] _1915_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__nand2_1
X_4760_ u_muldiv.o_div\[5\] _2173_ u_muldiv.o_div\[6\] vssd1 vssd1 vccd1 vccd1 _2178_
+ sky130_fd_sc_hd__o21ai_1
X_4691_ u_muldiv.divisor\[26\] u_muldiv.dividend\[26\] vssd1 vssd1 vccd1 vccd1 _2114_
+ sky130_fd_sc_hd__and2b_1
X_3711_ u_muldiv.mul\[41\] _1325_ _1438_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__a21oi_1
X_3642_ _1282_ _1288_ _1284_ _1281_ _0789_ _0920_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__mux4_1
X_5312_ u_muldiv.divisor\[24\] _2616_ _2617_ u_muldiv.divisor\[25\] vssd1 vssd1 vccd1
+ vccd1 _0415_ sky130_fd_sc_hd__a22o_1
X_3573_ _0653_ _0647_ _0650_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__mux2_1
X_5243_ _1029_ _2576_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__nand2_1
X_5174_ _2303_ _2510_ _2514_ vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__a21oi_1
X_4125_ _1711_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__clkbuf_4
X_4056_ u_bits.i_op2\[25\] u_bits.i_op2\[23\] _1681_ vssd1 vssd1 vccd1 vccd1 _1696_
+ sky130_fd_sc_hd__mux2_1
X_3007_ _0691_ _0692_ u_bits.i_op1\[24\] u_bits.i_op1\[25\] _0658_ _0659_ vssd1 vssd1
+ vccd1 vccd1 _0818_ sky130_fd_sc_hd__mux4_1
X_4958_ u_muldiv.divisor\[3\] u_muldiv.dividend\[3\] vssd1 vssd1 vccd1 vccd1 _2317_
+ sky130_fd_sc_hd__or2b_1
X_4889_ u_muldiv.quotient_msk\[1\] _1210_ _2279_ u_muldiv.quotient_msk\[2\] vssd1
+ vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__a22o_1
X_3909_ _0785_ i_op1[8] _1599_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_11_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_26_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4812_ _2208_ _2217_ _2218_ _2219_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__a31o_1
X_5792_ clknet_leaf_38_i_clk _0434_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[40\] sky130_fd_sc_hd__dfxtp_1
X_4743_ _2154_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__clkbuf_4
X_4674_ _2086_ _2096_ _2094_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__or3_1
X_3625_ _1106_ csr_data\[3\] _1124_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__o21ai_1
X_3556_ _0920_ _0948_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__nand2_1
X_5226_ _2556_ _2561_ _1877_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__mux2_1
X_3487_ o_wdata[1] _1233_ _0799_ u_wr_mux.i_reg_data2\[9\] vssd1 vssd1 vccd1 vccd1
+ _1235_ sky130_fd_sc_hd__a22o_1
X_5157_ _2036_ _2038_ _2098_ vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__and3_1
X_5088_ _2042_ _2043_ _2081_ vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__or3_1
X_4108_ u_pc_sel.i_pc_next\[14\] i_pc_next[14] _1723_ vssd1 vssd1 vccd1 vccd1 _1727_
+ sky130_fd_sc_hd__mux2_1
X_4039_ u_bits.i_op2\[20\] u_bits.i_op2\[18\] _1681_ vssd1 vssd1 vccd1 vccd1 _1684_
+ sky130_fd_sc_hd__mux2_1
X_3410_ _1141_ _1151_ _1180_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__and3_1
X_4390_ _1487_ _1852_ _1899_ _1856_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__a31o_1
X_3341_ _0528_ _0547_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__nor2_1
X_3272_ _0458_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__xnor2_1
X_5011_ _1880_ _2364_ _2365_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__and3_1
X_5775_ clknet_leaf_11_i_clk _0418_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_2987_ _0625_ _0799_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__and2_2
X_4726_ u_muldiv.divisor\[61\] u_muldiv.divisor\[60\] u_muldiv.divisor\[62\] u_muldiv.i_on_end
+ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__or4_1
X_4657_ u_muldiv.divisor\[13\] u_muldiv.dividend\[13\] vssd1 vssd1 vccd1 vccd1 _2080_
+ sky130_fd_sc_hd__or2b_1
X_3608_ _1337_ _1339_ _1340_ _1341_ _0789_ _0674_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__mux4_1
X_4588_ _2017_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__clkbuf_1
X_3539_ _1274_ o_add[0] _0804_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__a21oi_1
X_5209_ _2126_ u_muldiv.dividend\[24\] _2540_ _2111_ vssd1 vssd1 vccd1 vccd1 _2546_
+ sky130_fd_sc_hd__a22o_1
X_2910_ u_muldiv.dividend\[20\] _0721_ _0723_ u_muldiv.o_div\[20\] _0724_ vssd1 vssd1
+ vccd1 vccd1 _0725_ sky130_fd_sc_hd__a221o_1
X_3890_ _1594_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__buf_4
X_2841_ u_bits.i_op2\[0\] vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__clkbuf_4
X_5560_ clknet_leaf_7_i_clk _0207_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_2772_ _0456_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__xnor2_4
X_4511_ u_muldiv.mul\[15\] u_muldiv.mul\[16\] _1978_ vssd1 vssd1 vccd1 vccd1 _1987_
+ sky130_fd_sc_hd__mux2_1
X_5491_ clknet_leaf_51_i_clk _0139_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[9\]
+ sky130_fd_sc_hd__dfxtp_4
X_4442_ u_bits.i_op2\[22\] u_bits.i_op2\[23\] _1934_ vssd1 vssd1 vccd1 vccd1 _1942_
+ sky130_fd_sc_hd__or3_1
X_4373_ _1842_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__buf_2
X_3324_ _0702_ u_bits.i_op2\[31\] _0636_ _1116_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__o22a_1
X_3255_ _0644_ _1051_ _0712_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__o21a_1
X_3186_ u_bits.i_op1\[27\] u_muldiv.add_prev\[27\] _0451_ vssd1 vssd1 vccd1 vccd1
+ _0988_ sky130_fd_sc_hd__mux2_1
X_5758_ clknet_leaf_19_i_clk _0401_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4709_ u_muldiv.divisor\[29\] u_muldiv.dividend\[29\] vssd1 vssd1 vccd1 vccd1 _2132_
+ sky130_fd_sc_hd__or2b_1
X_5689_ clknet_leaf_26_i_clk _0332_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3040_ u_bits.i_op1\[23\] u_muldiv.add_prev\[23\] _0451_ vssd1 vssd1 vccd1 vccd1
+ _0850_ sky130_fd_sc_hd__mux2_1
X_4991_ _2056_ _2072_ _2071_ vssd1 vssd1 vccd1 vccd1 _2347_ sky130_fd_sc_hd__o21a_1
X_3942_ _1623_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__clkbuf_1
X_3873_ o_add[25] _1579_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__and2_1
X_5612_ clknet_leaf_34_i_clk _0259_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[29\] sky130_fd_sc_hd__dfxtp_1
X_2824_ _0638_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__clkbuf_2
X_5543_ clknet_leaf_16_i_clk _0191_ vssd1 vssd1 vccd1 vccd1 csr_data\[27\] sky130_fd_sc_hd__dfxtp_1
X_2755_ _0559_ _0560_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__nand2_1
X_2686_ u_bits.i_op1\[15\] u_muldiv.add_prev\[15\] _0449_ vssd1 vssd1 vccd1 vccd1
+ _0501_ sky130_fd_sc_hd__mux2_1
X_5474_ clknet_leaf_5_i_clk _0122_ vssd1 vssd1 vccd1 vccd1 o_funct3[0] sky130_fd_sc_hd__dfxtp_4
X_4425_ u_bits.i_op2\[20\] _1928_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__xnor2_1
X_4356_ u_bits.i_op2\[4\] _1376_ u_bits.i_op2\[6\] _1859_ vssd1 vssd1 vccd1 vccd1
+ _1873_ sky130_fd_sc_hd__or4_1
X_3307_ _1095_ _1100_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__nand2_1
X_4287_ _1818_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
X_3238_ _0858_ _1028_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__or3_1
X_3169_ _0644_ _0971_ _0712_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__o21a_1
X_4210_ u_wr_mux.i_reg_data2\[22\] i_reg_data2[22] _1778_ vssd1 vssd1 vccd1 vccd1
+ _1779_ sky130_fd_sc_hd__mux2_1
X_5190_ _2121_ _2528_ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__and2_1
X_4141_ _1742_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__clkbuf_1
X_4072_ u_bits.i_op2\[29\] _1687_ _1596_ i_op2[29] vssd1 vssd1 vccd1 vccd1 _1707_
+ sky130_fd_sc_hd__a22o_1
X_3023_ _0655_ u_bits.i_op1\[13\] _0658_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__mux2_1
X_4974_ u_muldiv.dividend\[4\] _2315_ vssd1 vssd1 vccd1 vccd1 _2332_ sky130_fd_sc_hd__xor2_1
X_3925_ _1614_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__clkbuf_1
X_3856_ _0672_ _1572_ _1573_ _0800_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__o211a_1
X_3787_ _1331_ _1506_ _1508_ _1509_ _0728_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__o221a_1
X_2807_ _0618_ _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__nor2_4
X_5526_ clknet_leaf_15_i_clk _0174_ vssd1 vssd1 vccd1 vccd1 csr_data\[10\] sky130_fd_sc_hd__dfxtp_1
X_2738_ _0448_ u_bits.i_op1\[7\] _0497_ _0552_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a31o_1
X_5457_ clknet_leaf_8_i_clk _0105_ vssd1 vssd1 vccd1 vccd1 o_res_src[1] sky130_fd_sc_hd__dfxtp_2
X_2669_ _0480_ _0483_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__nand2_1
X_4408_ u_bits.i_op2\[16\] _1910_ _1846_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__o21ai_1
X_5388_ clknet_leaf_49_i_clk _0036_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[20\] sky130_fd_sc_hd__dfxtp_2
X_4339_ u_bits.i_op2\[3\] _0916_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__or2_1
X_3710_ u_muldiv.dividend\[9\] _1326_ _1327_ u_muldiv.o_div\[9\] _1383_ vssd1 vssd1
+ vccd1 vccd1 _1438_ sky130_fd_sc_hd__a221o_1
X_4690_ u_muldiv.divisor\[27\] u_muldiv.dividend\[27\] vssd1 vssd1 vccd1 vccd1 _2113_
+ sky130_fd_sc_hd__xnor2_1
X_3641_ _1372_ _1373_ _1336_ u_pc_sel.i_pc_next\[4\] vssd1 vssd1 vccd1 vccd1 o_result[4]
+ sky130_fd_sc_hd__a2bb2o_2
X_3572_ u_bits.i_op1\[14\] u_bits.i_op1\[15\] _0650_ vssd1 vssd1 vccd1 vccd1 _1307_
+ sky130_fd_sc_hd__mux2_1
X_5311_ u_muldiv.divisor\[23\] _2616_ _2617_ u_muldiv.divisor\[24\] vssd1 vssd1 vccd1
+ vccd1 _0414_ sky130_fd_sc_hd__a22o_1
X_5242_ _0996_ _2568_ _2385_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__o21ai_1
X_5173_ _1206_ _2512_ _2513_ _1828_ vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__o31a_1
X_4124_ _1733_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__clkbuf_1
X_4055_ _1689_ _1694_ _1695_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__a21o_1
X_3006_ u_muldiv.mul\[22\] _0740_ _0741_ u_muldiv.mul\[54\] _0816_ vssd1 vssd1 vccd1
+ vccd1 _0817_ sky130_fd_sc_hd__a221o_1
X_4957_ u_muldiv.dividend\[3\] _2301_ vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__nand2_1
X_4888_ _1210_ u_muldiv.quotient_msk\[0\] _2279_ u_muldiv.quotient_msk\[1\] vssd1
+ vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__a22o_1
X_3908_ _1605_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__clkbuf_1
X_3839_ u_bits.i_op2\[18\] _0645_ _0637_ _1557_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__o22a_1
X_5509_ clknet_leaf_50_i_clk _0157_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[27\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_7_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4811_ u_muldiv.quotient_msk\[16\] u_muldiv.o_div\[16\] _1840_ vssd1 vssd1 vccd1
+ vccd1 _2219_ sky130_fd_sc_hd__o21a_1
X_5791_ clknet_leaf_38_i_clk _0433_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[39\] sky130_fd_sc_hd__dfxtp_1
X_4742_ _2157_ _2160_ _2163_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__o21a_1
X_4673_ _2087_ _2091_ _2090_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__a21o_1
X_3624_ _0454_ _1353_ _1355_ _1356_ _1357_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__o221a_1
X_3555_ _1285_ _1290_ _0687_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__mux2_1
X_3486_ _1192_ u_wr_mux.i_reg_data2\[24\] _1234_ vssd1 vssd1 vccd1 vccd1 o_wdata[24]
+ sky130_fd_sc_hd__a21o_2
X_5225_ _2558_ _2560_ _2288_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__mux2_1
X_5156_ u_muldiv.dividend\[20\] _2487_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__xor2_1
X_5087_ u_muldiv.dividend\[14\] _2423_ vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__xor2_1
X_4107_ _1726_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__clkbuf_1
X_4038_ _1665_ _1682_ _1683_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__a21o_1
X_3340_ _1130_ vssd1 vssd1 vccd1 vccd1 o_add[2] sky130_fd_sc_hd__inv_2
X_5010_ _2362_ _2363_ _1258_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__a21o_1
X_3271_ _0724_ u_bits.i_op2\[30\] _0465_ u_bits.i_op1\[30\] vssd1 vssd1 vccd1 vccd1
+ _1067_ sky130_fd_sc_hd__a22o_1
X_5774_ clknet_leaf_12_i_clk _0417_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_2986_ _0682_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__clkbuf_4
X_4725_ u_muldiv.divisor\[51\] u_muldiv.divisor\[50\] u_muldiv.divisor\[49\] u_muldiv.divisor\[48\]
+ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__or4_1
X_4656_ _2050_ _2051_ _2077_ _2048_ _2078_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__o311a_1
X_3607_ _1258_ _0785_ _1250_ _1305_ _0651_ _0774_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__mux4_1
X_4587_ o_add[31] _1584_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__and2_1
X_3538_ _1247_ _1264_ _1271_ _1273_ _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__a311o_1
X_3469_ _1225_ vssd1 vssd1 vccd1 vccd1 o_wdata[16] sky130_fd_sc_hd__buf_2
X_5208_ _2545_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__clkbuf_1
X_5139_ _2478_ _2480_ _2482_ _2288_ vssd1 vssd1 vccd1 vccd1 _2483_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_10_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_25_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2840_ u_bits.i_op1\[14\] vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__buf_4
X_2771_ _0449_ u_bits.i_op1\[10\] _0497_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__a31o_1
X_4510_ _1986_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__clkbuf_1
X_5490_ clknet_leaf_51_i_clk _0138_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[8\]
+ sky130_fd_sc_hd__dfxtp_4
X_4441_ u_muldiv.divisor\[54\] _1836_ _1887_ u_muldiv.divisor\[55\] _1941_ vssd1 vssd1
+ vccd1 vccd1 _0220_ sky130_fd_sc_hd__a221o_1
X_4372_ u_muldiv.divisor\[40\] _1867_ _1843_ u_muldiv.divisor\[41\] _1886_ vssd1 vssd1
+ vccd1 vccd1 _0206_ sky130_fd_sc_hd__a221o_1
X_3323_ _0617_ _0638_ _1115_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__and3_1
X_3254_ _0670_ _0765_ _0911_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__o21a_1
X_3185_ _0458_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__xnor2_1
X_5757_ clknet_leaf_26_i_clk _0400_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2969_ u_bits.i_op1\[15\] u_bits.i_op1\[14\] _0656_ vssd1 vssd1 vccd1 vccd1 _0782_
+ sky130_fd_sc_hd__mux2_1
X_4708_ _2122_ _2125_ _2129_ _2130_ _2030_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__o311ai_4
X_5688_ clknet_leaf_27_i_clk _0331_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4639_ u_muldiv.divisor\[1\] u_muldiv.dividend\[1\] vssd1 vssd1 vccd1 vccd1 _2062_
+ sky130_fd_sc_hd__xnor2_1
X_4990_ u_muldiv.dividend\[6\] _2336_ vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__nand2_1
X_3941_ _0692_ i_op1[23] _1621_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__mux2_1
X_3872_ _0903_ _1585_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__nor2_1
X_5611_ clknet_leaf_34_i_clk _0258_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[28\] sky130_fd_sc_hd__dfxtp_1
X_2823_ o_funct3[1] o_funct3[0] vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__nor2_2
X_5542_ clknet_leaf_16_i_clk _0190_ vssd1 vssd1 vccd1 vccd1 csr_data\[26\] sky130_fd_sc_hd__dfxtp_1
X_2754_ _0554_ _0555_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__nor2_1
X_5473_ clknet_leaf_14_i_clk _0121_ vssd1 vssd1 vccd1 vccd1 o_pc_target[15] sky130_fd_sc_hd__dfxtp_2
X_2685_ _0456_ _0499_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__xnor2_1
X_4424_ _1850_ _1927_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__nand2_1
X_4355_ u_muldiv.divisor\[37\] _1867_ _1843_ u_muldiv.divisor\[38\] _1872_ vssd1 vssd1
+ vccd1 vccd1 _0203_ sky130_fd_sc_hd__a221o_1
X_3306_ _0539_ _1099_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__xnor2_1
X_4286_ csr_data\[25\] i_csr_data[25] _1811_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__mux2_1
X_3237_ _0925_ _1031_ _1033_ _0914_ _1035_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__a221o_1
X_3168_ _0670_ _0970_ _0911_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__o21a_1
X_3099_ _0634_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__clkbuf_4
X_4140_ o_pc_target[13] i_pc_target[13] _1734_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__mux2_1
X_4071_ u_bits.i_op2\[30\] u_bits.i_op2\[28\] _1198_ vssd1 vssd1 vccd1 vccd1 _1706_
+ sky130_fd_sc_hd__mux2_1
X_3022_ _0645_ _0647_ _0653_ _0654_ _0651_ _0774_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__mux4_1
X_4973_ _1826_ _2326_ _2327_ _2329_ _2330_ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__a32o_1
X_3924_ _0654_ i_op1[15] _1610_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__mux2_1
X_3855_ _0687_ _1347_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__nand2_1
X_3786_ u_muldiv.mul\[14\] _0748_ _1400_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__o21ai_1
X_2806_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__or2_2
X_5525_ clknet_leaf_13_i_clk _0173_ vssd1 vssd1 vccd1 vccd1 csr_data\[9\] sky130_fd_sc_hd__dfxtp_1
X_2737_ u_mux.i_group_mux u_bits.i_op2\[7\] vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__and2b_1
X_5456_ clknet_leaf_51_i_clk _0104_ vssd1 vssd1 vccd1 vccd1 o_res_src[0] sky130_fd_sc_hd__dfxtp_2
X_2668_ _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__clkinv_2
X_4407_ u_muldiv.divisor\[47\] _1878_ _1829_ u_muldiv.divisor\[48\] _1914_ vssd1 vssd1
+ vccd1 vccd1 _0213_ sky130_fd_sc_hd__o221a_1
X_5387_ clknet_leaf_48_i_clk _0035_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[19\] sky130_fd_sc_hd__dfxtp_2
X_4338_ u_muldiv.divisor\[34\] _1838_ _1843_ u_muldiv.divisor\[35\] _1858_ vssd1 vssd1
+ vccd1 vccd1 _0200_ sky130_fd_sc_hd__a221o_1
X_4269_ csr_data\[17\] i_csr_data[17] _1800_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__mux2_1
X_3640_ _1106_ csr_data\[4\] _1124_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__o21ai_1
X_3571_ _1305_ _1251_ _0777_ _0776_ _0778_ _0783_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__mux4_1
X_5310_ u_muldiv.divisor\[22\] _2616_ _2617_ u_muldiv.divisor\[23\] vssd1 vssd1 vccd1
+ vccd1 _0413_ sky130_fd_sc_hd__a22o_1
X_5241_ _2303_ _2131_ _2574_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__nand3_1
X_5172_ _2295_ _2511_ _0768_ vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__a21oi_1
X_4123_ o_pc_target[5] i_pc_target[5] _1723_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__mux2_1
X_4054_ u_bits.i_op2\[23\] _1687_ _1675_ i_op2[23] vssd1 vssd1 vccd1 vccd1 _1695_
+ sky130_fd_sc_hd__a22o_1
X_3005_ u_muldiv.dividend\[22\] _0742_ _0743_ u_muldiv.o_div\[22\] _0744_ vssd1 vssd1
+ vccd1 vccd1 _0816_ sky130_fd_sc_hd__a221o_1
X_4956_ u_muldiv.dividend\[3\] _2301_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__or2_1
X_4887_ _1946_ vssd1 vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__buf_2
X_3907_ _1258_ i_op1[7] _1599_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__mux2_1
X_3838_ _0617_ _0639_ _1556_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__and3_1
X_5508_ clknet_leaf_50_i_clk _0156_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[26\]
+ sky130_fd_sc_hd__dfxtp_2
X_3769_ _0714_ _1491_ _1492_ _0623_ _1155_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__o32a_1
X_5439_ clknet_leaf_0_i_clk _0087_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[30\] sky130_fd_sc_hd__dfxtp_4
X_4810_ u_muldiv.o_div\[15\] u_muldiv.o_div\[16\] _2210_ vssd1 vssd1 vccd1 vccd1 _2218_
+ sky130_fd_sc_hd__or3_2
X_5790_ clknet_leaf_38_i_clk _0432_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[38\] sky130_fd_sc_hd__dfxtp_1
X_4741_ _2161_ _2162_ u_muldiv.o_div\[2\] vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__a21o_1
X_4672_ _2086_ _2093_ _2094_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__or3_1
X_3623_ _0728_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__buf_2
X_3554_ _0940_ _1289_ _0673_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__mux2_1
X_3485_ o_wdata[0] _1233_ _0799_ u_wr_mux.i_reg_data2\[8\] vssd1 vssd1 vccd1 vccd1
+ _1234_ sky130_fd_sc_hd__a22o_1
X_5224_ _0689_ _2559_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__xnor2_1
X_5155_ _2497_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__clkbuf_1
X_5086_ _2434_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__clkbuf_1
X_4106_ u_pc_sel.i_pc_next\[13\] i_pc_next[13] _1723_ vssd1 vssd1 vccd1 vccd1 _1726_
+ sky130_fd_sc_hd__mux2_1
X_4037_ u_bits.i_op2\[18\] _1663_ _1675_ i_op2[18] vssd1 vssd1 vccd1 vccd1 _1683_
+ sky130_fd_sc_hd__a22o_1
X_4939_ u_muldiv.dividend\[1\] _2299_ _2244_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__mux2_1
X_3270_ _0739_ csr_data\[29\] _1066_ _0732_ vssd1 vssd1 vccd1 vccd1 o_result[29] sky130_fd_sc_hd__o211a_2
X_5773_ clknet_leaf_12_i_clk _0416_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_4724_ u_muldiv.divisor\[59\] u_muldiv.divisor\[58\] u_muldiv.divisor\[57\] u_muldiv.divisor\[56\]
+ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__or4_1
X_2985_ _0672_ _0797_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__nand2_1
X_4655_ u_muldiv.divisor\[11\] u_muldiv.dividend\[11\] vssd1 vssd1 vccd1 vccd1 _2078_
+ sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_6_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3606_ _0794_ _1310_ _1257_ _0786_ _0651_ _0774_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__mux4_1
X_4586_ _2016_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__clkbuf_1
X_3537_ u_mux.i_add_override vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__buf_2
X_3468_ o_wdata[0] u_wr_mux.i_reg_data2\[16\] _1224_ vssd1 vssd1 vccd1 vccd1 _1225_
+ sky130_fd_sc_hd__mux2_1
X_5207_ u_muldiv.dividend\[24\] _2544_ _2485_ vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__mux2_1
X_3399_ _0523_ _0601_ _0608_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__nand3_2
X_5138_ _0645_ _2481_ vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__xnor2_1
X_5069_ _0777_ _2417_ _1839_ vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__o21a_1
X_2770_ u_mux.i_group_mux u_bits.i_op2\[10\] vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__and2b_1
X_4440_ _1939_ _1940_ _1833_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__a21oi_1
X_4371_ _1884_ _1885_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__nor2_1
X_3322_ _0702_ u_bits.i_op2\[31\] vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__nand2_1
X_3253_ u_muldiv.mul\[29\] _0740_ _0720_ u_muldiv.mul\[61\] _1049_ vssd1 vssd1 vccd1
+ vccd1 _1050_ sky130_fd_sc_hd__a221o_1
X_3184_ _0461_ u_bits.i_op2\[27\] _0465_ u_bits.i_op1\[27\] vssd1 vssd1 vccd1 vccd1
+ _0986_ sky130_fd_sc_hd__a22o_1
X_5756_ clknet_leaf_26_i_clk _0399_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_2968_ u_bits.i_op1\[17\] u_bits.i_op1\[16\] _0656_ vssd1 vssd1 vccd1 vccd1 _0781_
+ sky130_fd_sc_hd__mux2_1
X_5687_ clknet_leaf_28_i_clk _0330_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4707_ u_muldiv.dividend\[28\] u_muldiv.divisor\[28\] vssd1 vssd1 vccd1 vccd1 _2130_
+ sky130_fd_sc_hd__or2b_1
X_4638_ _2060_ u_muldiv.dividend\[2\] vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__or2_1
X_2899_ u_mux.i_add_override vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__buf_2
X_4569_ _2010_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__clkbuf_1
X_3940_ _1622_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__clkbuf_1
X_3871_ _0855_ _1585_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__nor2_1
X_5610_ clknet_leaf_33_i_clk _0257_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[27\] sky130_fd_sc_hd__dfxtp_1
X_2822_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__buf_2
X_5541_ clknet_leaf_15_i_clk _0189_ vssd1 vssd1 vccd1 vccd1 csr_data\[25\] sky130_fd_sc_hd__dfxtp_2
X_2753_ _0528_ _0547_ _0567_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__or3_2
X_5472_ clknet_leaf_14_i_clk _0120_ vssd1 vssd1 vccd1 vccd1 o_pc_target[14] sky130_fd_sc_hd__dfxtp_2
X_2684_ _0448_ u_bits.i_op1\[15\] _0497_ _0498_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__a31o_1
X_4423_ u_bits.i_op2\[18\] u_bits.i_op2\[19\] _1919_ vssd1 vssd1 vccd1 vccd1 _1927_
+ sky130_fd_sc_hd__or3_1
X_4354_ _1870_ _1871_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__nor2_1
X_3305_ _0452_ u_bits.i_op2\[31\] _1098_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__o21ai_1
X_4285_ _1817_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
X_3236_ _1029_ u_bits.i_op2\[28\] _0636_ _1034_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__o22a_1
X_3167_ _0822_ _0823_ _0668_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_24_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3098_ u_bits.i_op2\[24\] vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_39_i_clk clknet_2_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5739_ clknet_leaf_21_i_clk _0382_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[23\]
+ sky130_fd_sc_hd__dfxtp_2
X_4070_ _1689_ _1704_ _1705_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__a21o_1
X_3021_ _0691_ _0630_ _0768_ _0646_ _0779_ _0831_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__mux4_1
X_4972_ _1310_ _2295_ _2328_ _1826_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__a31oi_1
X_3923_ _1613_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__clkbuf_1
X_3854_ _0872_ _0876_ _0875_ _0880_ _0524_ _0789_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__mux4_1
X_2805_ o_funct3[0] vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__buf_4
X_3785_ u_muldiv.mul\[46\] _0741_ _1507_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__a21oi_1
X_5524_ clknet_leaf_12_i_clk _0172_ vssd1 vssd1 vccd1 vccd1 csr_data\[8\] sky130_fd_sc_hd__dfxtp_1
X_2736_ _0549_ _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__xnor2_1
X_5455_ clknet_leaf_10_i_clk _0103_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_2667_ _0478_ _0481_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__nand2_1
X_4406_ _1911_ _1912_ _1913_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__o21ai_1
X_5386_ clknet_leaf_48_i_clk _0034_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[18\] sky130_fd_sc_hd__dfxtp_2
X_4337_ _1855_ _1857_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__nor2_1
X_4268_ _1808_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__clkbuf_1
X_3219_ _0458_ _1018_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__xnor2_1
X_4199_ u_wr_mux.i_reg_data2\[17\] i_reg_data2[17] _1767_ vssd1 vssd1 vccd1 vccd1
+ _1773_ sky130_fd_sc_hd__mux2_1
X_3570_ u_bits.i_op1\[10\] vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__clkbuf_4
X_5240_ _2030_ _2130_ _2122_ _2125_ _2129_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__a2111o_1
X_5171_ _0768_ _2385_ _2511_ vssd1 vssd1 vccd1 vccd1 _2512_ sky130_fd_sc_hd__and3_1
X_4122_ _1732_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__clkbuf_1
X_4053_ _0905_ u_bits.i_op2\[22\] _1681_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__mux2_1
X_3004_ _0812_ _0815_ vssd1 vssd1 vccd1 vccd1 o_add[22] sky130_fd_sc_hd__xor2_4
X_4955_ _2314_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__clkbuf_1
X_3906_ _1604_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__clkbuf_1
X_4886_ _2167_ _2276_ _2278_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__a21oi_1
X_3837_ u_bits.i_op2\[18\] _0645_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__nand2_1
X_3768_ _1487_ _0776_ _0906_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__a21oi_2
X_5507_ clknet_leaf_50_i_clk _0155_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[25\]
+ sky130_fd_sc_hd__dfxtp_2
X_2719_ u_mux.i_group_mux _0533_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__and2b_1
X_3699_ _0454_ _1424_ _1426_ _1427_ _1357_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__o221a_1
X_5438_ clknet_leaf_0_i_clk _0086_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[29\] sky130_fd_sc_hd__dfxtp_4
X_5369_ clknet_leaf_47_i_clk _0017_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[1\] sky130_fd_sc_hd__dfxtp_1
X_4740_ _1835_ _2158_ u_muldiv.quotient_msk\[2\] vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__a21o_1
X_4671_ _2037_ _2036_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__or2b_1
X_3622_ u_muldiv.mul\[3\] _1330_ _1331_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__o21ai_1
X_3553_ _1288_ _0754_ _0696_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__mux2_1
X_3484_ _0718_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__buf_4
X_5223_ _0943_ _2548_ _2385_ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__o21ai_1
X_5154_ u_muldiv.dividend\[19\] _2496_ _2485_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__mux2_1
X_4105_ _1725_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__clkbuf_1
X_5085_ u_muldiv.dividend\[13\] _2433_ _2378_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__mux2_1
X_4036_ u_bits.i_op2\[19\] u_bits.i_op2\[17\] _1681_ vssd1 vssd1 vccd1 vccd1 _1682_
+ sky130_fd_sc_hd__mux2_1
X_4938_ _2208_ _2286_ _2287_ _2298_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__a31o_1
X_4869_ u_muldiv.quotient_msk\[28\] u_muldiv.o_div\[28\] _1840_ vssd1 vssd1 vccd1
+ vccd1 _2265_ sky130_fd_sc_hd__o21a_1
X_5772_ clknet_leaf_11_i_clk _0415_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_2984_ _0669_ _0793_ _0796_ _0707_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__a211o_1
X_4723_ u_muldiv.divisor\[40\] _2140_ _2145_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__or3_1
X_4654_ _2054_ _2055_ _2075_ _2052_ _2076_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__o311a_1
X_3605_ _1338_ _1286_ _0779_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__mux2_1
X_4585_ o_add[30] _2004_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__and2_1
X_3536_ _0831_ _0917_ _1272_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__a21oi_1
X_5206_ _2536_ _2543_ _1877_ vssd1 vssd1 vccd1 vccd1 _2544_ sky130_fd_sc_hd__mux2_1
X_3467_ _0619_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__buf_4
X_3398_ o_add[11] o_add[14] o_add[18] vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__or3_1
X_5137_ _0647_ _2469_ _2385_ vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__o21ai_1
X_5068_ _0777_ _2417_ vssd1 vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__nand2_1
X_4019_ u_bits.i_op2\[14\] u_bits.i_op2\[12\] _1657_ vssd1 vssd1 vccd1 vccd1 _1670_
+ sky130_fd_sc_hd__mux2_1
X_4370_ u_bits.i_op2\[9\] _1852_ _1883_ _1856_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__a31o_1
X_3321_ _0873_ _1113_ _0674_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__mux2_1
X_3252_ u_muldiv.dividend\[29\] _0721_ _0723_ u_muldiv.o_div\[29\] _0744_ vssd1 vssd1
+ vccd1 vccd1 _1049_ sky130_fd_sc_hd__a221o_1
X_3183_ _0739_ csr_data\[26\] _0985_ _0732_ vssd1 vssd1 vccd1 vccd1 o_result[26] sky130_fd_sc_hd__o211a_2
X_5755_ clknet_leaf_26_i_clk _0398_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2967_ _0776_ _0777_ u_bits.i_op1\[11\] u_bits.i_op1\[10\] _0778_ _0779_ vssd1 vssd1
+ vccd1 vccd1 _0780_ sky130_fd_sc_hd__mux4_2
X_5686_ clknet_leaf_28_i_clk _0329_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4706_ _2118_ _2128_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__nor2_1
X_2898_ _0688_ _0709_ _0712_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__o21ai_1
X_4637_ u_muldiv.divisor\[2\] vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__inv_2
X_4568_ o_add[19] _2004_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__and2_1
X_4499_ u_muldiv.mul\[9\] u_muldiv.mul\[10\] _1978_ vssd1 vssd1 vccd1 vccd1 _1981_
+ sky130_fd_sc_hd__mux2_1
X_3519_ _0917_ _0791_ _1255_ _0794_ _0831_ _1112_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_5_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3870_ _1584_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__clkbuf_4
X_2821_ _0620_ _0635_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__nor2_4
X_5540_ clknet_leaf_15_i_clk _0188_ vssd1 vssd1 vccd1 vccd1 csr_data\[24\] sky130_fd_sc_hd__dfxtp_1
X_2752_ _0551_ _0562_ _0566_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__or3_1
X_5471_ clknet_leaf_14_i_clk _0119_ vssd1 vssd1 vccd1 vccd1 o_pc_target[13] sky130_fd_sc_hd__dfxtp_2
X_2683_ u_mux.i_group_mux u_bits.i_op2\[15\] vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__and2b_1
X_4422_ u_muldiv.divisor\[50\] _1836_ _1887_ u_muldiv.divisor\[51\] _1926_ vssd1 vssd1
+ vccd1 vccd1 _0216_ sky130_fd_sc_hd__a221o_1
X_4353_ u_bits.i_op2\[6\] _1850_ _1869_ _1856_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__a31o_1
X_4284_ csr_data\[24\] i_csr_data[24] _1811_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__mux2_1
X_3304_ _1096_ _1097_ _0452_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__o21ai_1
X_3235_ _1029_ u_bits.i_op2\[28\] _0867_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__a21oi_1
X_3166_ u_muldiv.mul\[26\] _0740_ _0741_ u_muldiv.mul\[58\] _0968_ vssd1 vssd1 vccd1
+ vccd1 _0969_ sky130_fd_sc_hd__a221o_1
X_3097_ u_bits.i_op1\[24\] vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__clkbuf_4
X_3999_ _1406_ _1637_ _1651_ i_op2[7] vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__a22o_1
X_5738_ clknet_leaf_21_i_clk _0381_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[22\]
+ sky130_fd_sc_hd__dfxtp_2
X_5669_ clknet_leaf_29_i_clk _0312_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[15\] sky130_fd_sc_hd__dfxtp_1
X_3020_ _0778_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__buf_4
X_4971_ _2295_ _2328_ _1310_ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__a21o_1
X_3922_ _0655_ i_op1[14] _1610_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__mux2_1
X_3853_ u_bits.i_op2\[19\] _0646_ _0637_ _1570_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__o22a_1
X_2804_ o_funct3[1] vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__buf_4
X_3784_ u_muldiv.dividend\[14\] _0742_ _0743_ u_muldiv.o_div\[14\] _1383_ vssd1 vssd1
+ vccd1 vccd1 _1507_ sky130_fd_sc_hd__a221o_1
X_5523_ clknet_leaf_12_i_clk _0171_ vssd1 vssd1 vccd1 vccd1 csr_data\[7\] sky130_fd_sc_hd__dfxtp_1
X_2735_ u_bits.i_op1\[4\] u_muldiv.add_prev\[4\] _0450_ vssd1 vssd1 vccd1 vccd1 _0550_
+ sky130_fd_sc_hd__mux2_1
X_5454_ clknet_leaf_10_i_clk _0102_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_2666_ _0476_ _0477_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__or2_1
X_5385_ clknet_leaf_48_i_clk _0033_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[17\] sky130_fd_sc_hd__dfxtp_2
X_4405_ _1880_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__buf_4
X_4336_ _0909_ _0916_ _1852_ _1856_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__a31o_1
X_4267_ csr_data\[16\] i_csr_data[16] _1800_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__mux2_1
X_4198_ _1772_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__clkbuf_1
X_3218_ _0461_ u_bits.i_op2\[28\] _0465_ u_bits.i_op1\[28\] vssd1 vssd1 vccd1 vccd1
+ _1018_ sky130_fd_sc_hd__a22o_1
X_3149_ _0628_ _0942_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_23_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5170_ u_bits.i_op1\[20\] u_bits.i_op1\[19\] _2492_ vssd1 vssd1 vccd1 vccd1 _2511_
+ sky130_fd_sc_hd__or3_2
X_4121_ o_pc_target[4] i_pc_target[4] _1723_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_i_clk clknet_2_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4052_ _1689_ _1692_ _1693_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__a21o_1
X_3003_ _0737_ _0736_ _0814_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__o21ai_2
X_4954_ u_muldiv.dividend\[2\] _2313_ _2244_ vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__mux2_1
X_3905_ _0786_ i_op1[6] _1599_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__mux2_1
X_4885_ _2161_ _2277_ u_muldiv.o_div\[31\] vssd1 vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__a21oi_1
X_3836_ _0751_ _1316_ _0711_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__o21a_1
X_3767_ _0908_ _1490_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__nor2_1
X_5506_ clknet_leaf_50_i_clk _0154_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[24\]
+ sky130_fd_sc_hd__dfxtp_2
X_2718_ u_bits.i_op2\[1\] vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__clkbuf_4
X_3698_ u_muldiv.mul\[8\] _1330_ _1400_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__o21ai_1
X_2649_ _0463_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__buf_2
X_5437_ clknet_leaf_0_i_clk _0085_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[28\] sky130_fd_sc_hd__dfxtp_4
X_5368_ clknet_leaf_47_i_clk _0016_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[0\] sky130_fd_sc_hd__dfxtp_2
X_5299_ u_muldiv.divisor\[13\] _2614_ _2615_ u_muldiv.divisor\[14\] vssd1 vssd1 vccd1
+ vccd1 _0404_ sky130_fd_sc_hd__a22o_1
X_4319_ _1841_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__buf_4
X_4670_ _2089_ _2092_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__or2b_1
X_3621_ u_muldiv.mul\[35\] _1325_ _1354_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__a21oi_1
X_3552_ _1286_ _1287_ _0648_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__mux2_1
X_3483_ _1232_ vssd1 vssd1 vccd1 vccd1 o_wdata[23] sky130_fd_sc_hd__buf_2
X_5222_ _2116_ _2557_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__xnor2_1
X_5153_ _1208_ _2487_ _2488_ _2491_ _2495_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__a32o_1
X_4104_ u_pc_sel.i_pc_next\[12\] i_pc_next[12] _1723_ vssd1 vssd1 vccd1 vccd1 _1725_
+ sky130_fd_sc_hd__mux2_1
X_5084_ _1208_ _2423_ _2424_ _2432_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__a31o_1
X_4035_ _1198_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__clkbuf_4
X_4937_ _2229_ _2297_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__nor2_1
X_4868_ u_muldiv.o_div\[27\] u_muldiv.o_div\[28\] _2258_ vssd1 vssd1 vccd1 vccd1 _2264_
+ sky130_fd_sc_hd__or3_2
X_3819_ _1106_ csr_data\[16\] _1539_ _1124_ vssd1 vssd1 vccd1 vccd1 o_result[16] sky130_fd_sc_hd__o211a_2
X_4799_ u_muldiv.o_div\[13\] _2201_ u_muldiv.o_div\[14\] vssd1 vssd1 vccd1 vccd1 _2209_
+ sky130_fd_sc_hd__o21ai_1
X_5771_ clknet_leaf_12_i_clk _0414_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_2983_ _0668_ _0795_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__nor2_1
X_4722_ _2141_ _2142_ _2143_ _2144_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__or4_1
X_4653_ u_muldiv.divisor\[9\] u_muldiv.dividend\[9\] vssd1 vssd1 vccd1 vccd1 _2076_
+ sky130_fd_sc_hd__or2b_1
X_3604_ u_bits.i_op1\[15\] _0653_ _0650_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__mux2_1
X_4584_ _2015_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__clkbuf_1
X_3535_ _0634_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__buf_2
X_3466_ _1223_ vssd1 vssd1 vccd1 vccd1 o_wdata[15] sky130_fd_sc_hd__buf_2
X_5205_ _2303_ _2538_ _2539_ _2541_ _2542_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__o32ai_1
X_3397_ o_add[21] o_add[22] o_add[15] o_add[19] vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__or4_1
X_5136_ _1826_ _2479_ vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__nand2_1
X_5067_ _1305_ _1251_ _2394_ _2292_ vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__o31a_1
X_4018_ _1665_ _1668_ _1669_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__a21o_1
X_3320_ _1111_ _1056_ _1001_ _0944_ _1112_ _0825_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__mux4_1
X_3251_ _1047_ _1048_ vssd1 vssd1 vccd1 vccd1 o_add[29] sky130_fd_sc_hd__xnor2_4
X_3182_ _0969_ _0984_ _0447_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__a21o_1
X_5754_ clknet_leaf_26_i_clk _0397_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2966_ _0663_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__buf_4
X_4705_ _2108_ _2127_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__or2_1
X_5685_ clknet_leaf_36_i_clk _0328_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[31\] sky130_fd_sc_hd__dfxtp_1
X_2897_ _0711_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__buf_2
X_4636_ u_muldiv.dividend\[3\] u_muldiv.divisor\[3\] vssd1 vssd1 vccd1 vccd1 _2059_
+ sky130_fd_sc_hd__or2b_1
X_4567_ _2009_ _2007_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__nor2_1
X_4498_ _1980_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
X_3518_ u_bits.i_op1\[2\] vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__clkbuf_4
X_3449_ _1194_ _1213_ _1214_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__mux2_1
X_5119_ _2464_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__clkbuf_1
X_2820_ _0619_ o_funct3[2] vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__nand2_1
X_2751_ _0564_ _0565_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__xnor2_4
X_5470_ clknet_leaf_14_i_clk _0118_ vssd1 vssd1 vccd1 vccd1 o_pc_target[12] sky130_fd_sc_hd__dfxtp_2
X_2682_ _0462_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__buf_2
X_4421_ _1924_ _1925_ _1833_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__a21oi_1
X_4352_ _1868_ _1869_ u_bits.i_op2\[6\] vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__a21oi_1
X_4283_ _1816_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__clkbuf_1
X_3303_ u_bits.i_op1\[31\] _0497_ _0626_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__a21oi_1
X_3234_ _1032_ _0680_ _0524_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__mux2_1
X_3165_ u_muldiv.dividend\[26\] _0742_ _0743_ u_muldiv.o_div\[26\] _0744_ vssd1 vssd1
+ vccd1 vccd1 _0968_ sky130_fd_sc_hd__a221o_1
X_3096_ _0903_ vssd1 vssd1 vccd1 vccd1 o_add[24] sky130_fd_sc_hd__inv_2
X_3998_ u_bits.i_op2\[8\] u_bits.i_op2\[6\] _1639_ vssd1 vssd1 vccd1 vccd1 _1655_
+ sky130_fd_sc_hd__mux2_1
X_5737_ clknet_leaf_17_i_clk _0380_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[21\]
+ sky130_fd_sc_hd__dfxtp_2
X_2949_ _0663_ _0703_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__nand2_1
X_5668_ clknet_leaf_29_i_clk _0311_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[14\] sky130_fd_sc_hd__dfxtp_1
X_4619_ _2040_ _2041_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__nand2_1
X_5599_ clknet_leaf_35_i_clk _0246_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[16\] sky130_fd_sc_hd__dfxtp_1
X_4970_ u_bits.i_op1\[2\] u_bits.i_op1\[3\] _2308_ vssd1 vssd1 vccd1 vccd1 _2328_
+ sky130_fd_sc_hd__or3_4
X_3921_ _1612_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__clkbuf_1
X_3852_ _0617_ _0639_ _1569_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__and3_1
X_2803_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__clkbuf_4
X_5522_ clknet_leaf_12_i_clk _0170_ vssd1 vssd1 vccd1 vccd1 csr_data\[6\] sky130_fd_sc_hd__dfxtp_1
X_3783_ _0714_ _1504_ _1505_ _0623_ _1163_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__o32a_1
X_2734_ _0456_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__xnor2_1
X_5453_ clknet_leaf_10_i_clk _0101_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_2665_ _0479_ _0474_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__nor2_2
X_5384_ clknet_leaf_48_i_clk _0032_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[16\] sky130_fd_sc_hd__dfxtp_2
X_4404_ u_bits.i_op2\[16\] _1846_ _1910_ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__and3_1
X_4335_ _1831_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__buf_2
X_4266_ _1807_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__clkbuf_1
X_4197_ u_wr_mux.i_reg_data2\[16\] i_reg_data2[16] _1767_ vssd1 vssd1 vccd1 vccd1
+ _1772_ sky130_fd_sc_hd__mux2_1
X_3217_ _1015_ _1016_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__nand2_1
X_3148_ _0925_ _0946_ _0949_ _0914_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__a221o_1
X_3079_ _0750_ o_add[23] _0887_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_4_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4120_ _1731_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__clkbuf_1
X_4051_ u_bits.i_op2\[22\] _1687_ _1675_ i_op2[22] vssd1 vssd1 vccd1 vccd1 _1693_
+ sky130_fd_sc_hd__a22o_1
X_3002_ _0734_ _0735_ _0813_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o21ai_1
X_4953_ _2208_ _2301_ _2302_ _2312_ vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__a31o_1
X_3904_ _1603_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__clkbuf_1
X_4884_ u_muldiv.quotient_msk\[31\] _1878_ _2271_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__a21o_1
X_3835_ u_muldiv.mul\[18\] _0717_ _0720_ u_muldiv.mul\[50\] _1553_ vssd1 vssd1 vccd1
+ vccd1 _1554_ sky130_fd_sc_hd__a221o_1
X_3766_ _1110_ _1055_ _1486_ _1248_ _1489_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__a221o_1
X_2717_ _0530_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__xnor2_1
X_5505_ clknet_leaf_47_i_clk _0153_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[23\]
+ sky130_fd_sc_hd__dfxtp_2
X_3697_ u_muldiv.mul\[40\] _1325_ _1425_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__a21oi_1
X_5436_ clknet_leaf_1_i_clk _0084_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[27\] sky130_fd_sc_hd__dfxtp_4
X_2648_ u_mux.i_group_mux _0462_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__and2_1
X_5367_ clknet_leaf_23_i_clk _0015_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[63\] sky130_fd_sc_hd__dfxtp_1
X_5298_ u_muldiv.divisor\[12\] _2614_ _2615_ u_muldiv.divisor\[13\] vssd1 vssd1 vccd1
+ vccd1 _0403_ sky130_fd_sc_hd__a22o_1
X_4318_ _1840_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__buf_4
X_4249_ _1798_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
X_3620_ u_muldiv.dividend\[3\] _1326_ _1327_ u_muldiv.o_div\[3\] _0717_ vssd1 vssd1
+ vccd1 vccd1 _1354_ sky130_fd_sc_hd__a221o_1
X_3551_ u_bits.i_op1\[19\] _0630_ _0657_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__mux2_1
X_3482_ o_wdata[7] u_wr_mux.i_reg_data2\[23\] _1224_ vssd1 vssd1 vccd1 vccd1 _1232_
+ sky130_fd_sc_hd__mux2_1
X_5221_ _2120_ _2528_ _2112_ _2128_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__o31ai_2
X_5152_ _1827_ _2493_ _2494_ _1840_ vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__a31o_1
X_4103_ _1724_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__clkbuf_1
X_5083_ _2426_ _2427_ _2431_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__o21a_1
X_4034_ _1665_ _1679_ _1680_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__a21o_1
X_4936_ _2288_ _2289_ _2290_ _2294_ _2296_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__o32a_1
X_4867_ u_muldiv.o_div\[27\] _2258_ u_muldiv.o_div\[28\] vssd1 vssd1 vccd1 vccd1 _2263_
+ sky130_fd_sc_hd__o21ai_1
X_3818_ _1527_ _1538_ _0446_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__a21o_1
X_4798_ _1207_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__buf_4
X_3749_ u_bits.i_op2\[12\] _0777_ _1267_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__a21oi_1
X_5419_ clknet_leaf_49_i_clk _0067_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[10\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_22_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_37_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5770_ clknet_leaf_12_i_clk _0413_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_2982_ u_bits.i_op1\[5\] u_bits.i_op1\[4\] _0794_ u_bits.i_op1\[2\] _0650_ _0648_
+ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__mux4_2
X_4721_ _1834_ u_muldiv.dividend\[31\] vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__nor2_1
X_4652_ _2056_ _2071_ _2072_ _2074_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__o31a_1
X_3603_ _1251_ _0777_ _0776_ _0655_ _0778_ _0779_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__mux4_1
X_4583_ o_add[29] _2004_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__and2_1
X_3534_ _1265_ _1266_ _1270_ _0906_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__o211a_1
X_3465_ u_wr_mux.i_reg_data2\[15\] o_wdata[7] _0718_ vssd1 vssd1 vccd1 vccd1 _1223_
+ sky130_fd_sc_hd__mux2_1
X_5204_ _2540_ _2111_ _2303_ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__o21ai_1
X_3396_ u_adder.i_cmp_inverse vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__clkinv_2
X_5135_ _2096_ _2477_ _2086_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__a21o_1
X_5066_ _2047_ _2079_ _2046_ vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__o21ai_1
X_4017_ u_bits.i_op2\[12\] _1663_ _1651_ i_op2[12] vssd1 vssd1 vccd1 vccd1 _1669_
+ sky130_fd_sc_hd__a22o_1
X_4919_ _1209_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__clkbuf_4
X_3250_ _1017_ _1023_ _1021_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__a21bo_1
X_3181_ _0750_ o_add[26] _0982_ _0983_ _0804_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__a221o_1
X_5753_ clknet_leaf_25_i_clk _0396_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4704_ _2126_ u_muldiv.dividend\[24\] _2107_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__a21oi_1
X_2965_ _0657_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__buf_4
X_5684_ clknet_leaf_36_i_clk _0327_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[30\] sky130_fd_sc_hd__dfxtp_1
X_2896_ _0642_ _0703_ _0710_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__a21oi_4
X_4635_ u_muldiv.dividend\[4\] u_muldiv.divisor\[4\] vssd1 vssd1 vccd1 vccd1 _2058_
+ sky130_fd_sc_hd__or2b_1
X_4566_ o_add[18] vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__inv_2
X_3517_ _1252_ _1253_ _0760_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__mux2_1
X_4497_ u_muldiv.mul\[8\] u_muldiv.mul\[9\] _1978_ vssd1 vssd1 vccd1 vccd1 _1980_
+ sky130_fd_sc_hd__mux2_1
X_3448_ _1198_ u_muldiv.i_on_wait vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__nor2_8
X_3379_ _0505_ _0506_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__or2_1
X_5118_ u_muldiv.dividend\[16\] _2463_ _2378_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__mux2_1
X_5049_ _1878_ _2393_ _2400_ vssd1 vssd1 vccd1 vccd1 _2401_ sky130_fd_sc_hd__o21a_1
X_2750_ u_bits.i_op1\[5\] u_muldiv.add_prev\[5\] _0450_ vssd1 vssd1 vccd1 vccd1 _0565_
+ sky130_fd_sc_hd__mux2_2
X_2681_ _0474_ _0478_ _0484_ _0494_ _0495_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__o221a_1
X_4420_ u_bits.i_op2\[19\] _1923_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__or2_1
X_4351_ _0688_ _1376_ _1859_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__or3_1
X_4282_ csr_data\[23\] i_csr_data[23] _1811_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__mux2_1
X_3302_ u_bits.i_op1\[31\] _0497_ _0626_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__and3_1
X_3233_ _0664_ _0667_ _0696_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__mux2_1
X_3164_ _0964_ _0967_ vssd1 vssd1 vccd1 vccd1 o_add[26] sky130_fd_sc_hd__xor2_4
X_3095_ _0901_ _0902_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__nand2_1
X_3997_ _1641_ _1653_ _1654_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__a21o_1
X_5736_ clknet_leaf_16_i_clk _0379_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[20\]
+ sky130_fd_sc_hd__dfxtp_2
X_2948_ _0697_ _0699_ _0656_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__mux2_1
X_5667_ clknet_leaf_29_i_clk _0310_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[13\] sky130_fd_sc_hd__dfxtp_1
X_4618_ u_muldiv.dividend\[14\] u_muldiv.divisor\[14\] vssd1 vssd1 vccd1 vccd1 _2041_
+ sky130_fd_sc_hd__or2b_1
X_2879_ _0668_ _0693_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__and2b_1
X_5598_ clknet_leaf_35_i_clk _0245_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[15\] sky130_fd_sc_hd__dfxtp_1
X_4549_ _1128_ _2006_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__nor2_1
X_3920_ _0776_ i_op1[13] _1610_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__mux2_1
X_3851_ u_bits.i_op2\[19\] _0646_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__nand2_1
X_2802_ o_funct3[2] vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__clkbuf_4
X_3782_ u_bits.i_op2\[14\] _0655_ _0906_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__a21oi_1
X_5521_ clknet_leaf_12_i_clk _0169_ vssd1 vssd1 vccd1 vccd1 csr_data\[5\] sky130_fd_sc_hd__dfxtp_1
X_2733_ _0459_ u_bits.i_op2\[4\] u_bits.i_op1\[4\] _0463_ vssd1 vssd1 vccd1 vccd1
+ _0548_ sky130_fd_sc_hd__a22o_1
X_5452_ clknet_leaf_10_i_clk _0100_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_2664_ _0472_ _0473_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__and2_1
X_5383_ clknet_leaf_48_i_clk _0031_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[15\] sky130_fd_sc_hd__dfxtp_2
X_4403_ _1868_ _1910_ u_bits.i_op2\[16\] vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__a21oi_1
X_4334_ _0916_ _1850_ _0909_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__a21oi_1
X_4265_ csr_data\[15\] i_csr_data[15] _1800_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__mux2_1
X_4196_ _1771_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__clkbuf_1
X_3216_ _0895_ _0896_ _0900_ _0936_ _1013_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__a2111o_1
X_3147_ _0943_ u_bits.i_op2\[25\] _0636_ _0951_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__o22a_1
X_3078_ _0747_ _0885_ _0886_ _0453_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__a31o_1
X_5719_ clknet_leaf_24_i_clk _0362_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4050_ u_bits.i_op2\[23\] u_bits.i_op2\[21\] _1681_ vssd1 vssd1 vccd1 vccd1 _1692_
+ sky130_fd_sc_hd__mux2_1
X_3001_ _0467_ _0468_ _0734_ _0735_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__a22o_1
X_4952_ _2303_ _2307_ _2311_ vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__a21oi_1
X_4883_ u_muldiv.o_div\[31\] _2271_ _1913_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__a21o_1
X_3903_ _1257_ i_op1[5] _1599_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__mux2_1
X_3834_ u_muldiv.dividend\[18\] _0721_ _0723_ u_muldiv.o_div\[18\] _0724_ vssd1 vssd1
+ vccd1 vccd1 _1553_ sky130_fd_sc_hd__a221o_1
X_3765_ _1487_ _0776_ _0926_ _1488_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__o22a_1
X_3696_ u_muldiv.dividend\[8\] _1326_ _1327_ u_muldiv.o_div\[8\] _1383_ vssd1 vssd1
+ vccd1 vccd1 _1425_ sky130_fd_sc_hd__a221o_1
X_2716_ u_bits.i_op1\[2\] u_muldiv.add_prev\[2\] _0450_ vssd1 vssd1 vccd1 vccd1 _0531_
+ sky130_fd_sc_hd__mux2_1
X_5504_ clknet_leaf_47_i_clk _0152_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[22\]
+ sky130_fd_sc_hd__dfxtp_2
X_2647_ u_bits.i_op2\[0\] u_bits.i_op2\[31\] u_muldiv.i_is_div vssd1 vssd1 vccd1 vccd1
+ _0462_ sky130_fd_sc_hd__mux2_1
X_5435_ clknet_leaf_1_i_clk _0083_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[26\] sky130_fd_sc_hd__dfxtp_4
X_5366_ clknet_leaf_34_i_clk _0014_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[62\] sky130_fd_sc_hd__dfxtp_1
X_5297_ u_muldiv.divisor\[11\] _2614_ _2615_ u_muldiv.divisor\[12\] vssd1 vssd1 vccd1
+ vccd1 _0402_ sky130_fd_sc_hd__a22o_1
X_4317_ _1839_ _1206_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__nor2_8
X_4248_ csr_data\[7\] i_csr_data[7] _1789_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__mux2_1
X_4179_ _1762_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__clkbuf_1
X_3550_ u_bits.i_op1\[17\] _0645_ _0657_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__mux2_1
X_5220_ u_muldiv.dividend\[26\] _2552_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__xor2_1
X_3481_ _1231_ vssd1 vssd1 vccd1 vccd1 o_wdata[22] sky130_fd_sc_hd__buf_2
X_5151_ _2295_ _2492_ _0646_ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__a21o_1
X_5082_ _1827_ _2429_ _2430_ _1840_ vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__a31o_1
X_4102_ u_pc_sel.i_pc_next\[11\] i_pc_next[11] _1723_ vssd1 vssd1 vccd1 vccd1 _1724_
+ sky130_fd_sc_hd__mux2_1
X_4033_ u_bits.i_op2\[17\] _1663_ _1675_ i_op2[17] vssd1 vssd1 vccd1 vccd1 _1680_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_3_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4935_ _0917_ _2295_ _0791_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__a21oi_1
X_4866_ _2167_ _2260_ _2262_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__a21oi_1
X_4797_ _2181_ _2205_ _2207_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__a21oi_1
X_3817_ _0749_ o_add[16] _1536_ _1537_ _0453_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__a221o_1
X_3748_ _0687_ _1027_ _1471_ _1472_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__a22o_1
X_3679_ _0674_ _0925_ _0882_ _1408_ _0858_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__a311o_1
X_5418_ clknet_leaf_51_i_clk _0066_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[9\] sky130_fd_sc_hd__dfxtp_4
X_5349_ o_add[16] _1214_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__and2_1
X_2981_ u_bits.i_op1\[3\] vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__clkbuf_4
X_4720_ u_muldiv.divisor\[47\] u_muldiv.divisor\[46\] u_muldiv.divisor\[45\] u_muldiv.divisor\[44\]
+ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__or4_1
X_4651_ _2073_ _2056_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__nor2_1
X_3602_ _1334_ _1335_ _1336_ u_pc_sel.i_pc_next\[2\] vssd1 vssd1 vccd1 vccd1 o_result[2]
+ sky130_fd_sc_hd__a2bb2o_2
X_4582_ _1024_ _1579_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__nor2_1
X_3533_ _0622_ o_add[0] _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__a21oi_1
X_3464_ _1222_ vssd1 vssd1 vccd1 vccd1 o_wdata[14] sky130_fd_sc_hd__buf_2
X_5203_ _2540_ _2111_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__and2_1
X_5134_ _2086_ _2096_ _2477_ vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__and3_1
X_3395_ u_adder.i_cmp_inverse _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__xnor2_1
X_5065_ _2046_ _2047_ _2079_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__or3_1
X_4016_ _1487_ u_bits.i_op2\[11\] _1657_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__mux2_1
X_4918_ u_muldiv.quotient_msk\[26\] _2282_ _2283_ u_muldiv.quotient_msk\[27\] vssd1
+ vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__a22o_1
X_4849_ u_muldiv.o_div\[23\] _2241_ u_muldiv.o_div\[24\] vssd1 vssd1 vccd1 vccd1 _2249_
+ sky130_fd_sc_hd__o21ai_1
X_3180_ _0629_ _0978_ _0955_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__a21oi_1
X_5752_ clknet_leaf_25_i_clk _0395_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2964_ u_bits.i_op1\[12\] vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__buf_4
X_4703_ u_muldiv.divisor\[24\] vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__inv_2
X_5683_ clknet_leaf_32_i_clk _0326_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[29\] sky130_fd_sc_hd__dfxtp_1
X_2895_ _0617_ _0682_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__nand2_2
X_4634_ u_muldiv.dividend\[5\] u_muldiv.divisor\[5\] vssd1 vssd1 vccd1 vccd1 _2057_
+ sky130_fd_sc_hd__and2b_1
X_4565_ _1176_ _2007_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__nor2_1
X_3516_ u_bits.i_op1\[12\] u_bits.i_op1\[13\] _0655_ u_bits.i_op1\[15\] _0650_ _0648_
+ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_21_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4496_ _1979_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
X_3447_ i_funct3[0] i_funct3[1] vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__nand2_1
X_3378_ _0508_ _0502_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__or2_2
X_5117_ _2457_ _2462_ _1877_ vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__mux2_1
X_5048_ _2375_ _2395_ _2396_ _1207_ _2399_ vssd1 vssd1 vccd1 vccd1 _2400_ sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_36_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2680_ _0472_ _0473_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__nand2_1
X_4350_ _1846_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__buf_2
X_3301_ _0702_ u_muldiv.add_prev\[31\] _0452_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__mux2_1
X_4281_ _1815_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__clkbuf_1
X_3232_ _0652_ _0660_ _1030_ _0922_ _0668_ _0673_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__mux4_1
X_3163_ _0901_ _0936_ _0966_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__o21ai_4
X_3094_ _0895_ _0896_ _0900_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__nand3_1
X_3996_ u_bits.i_op2\[6\] _1637_ _1651_ i_op2[6] vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__a22o_1
X_5735_ clknet_leaf_18_i_clk _0378_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[19\]
+ sky130_fd_sc_hd__dfxtp_2
X_2947_ _0696_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__buf_4
X_5666_ clknet_leaf_29_i_clk _0309_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[12\] sky130_fd_sc_hd__dfxtp_1
X_4617_ u_muldiv.divisor\[14\] u_muldiv.dividend\[14\] vssd1 vssd1 vccd1 vccd1 _2040_
+ sky130_fd_sc_hd__or2b_1
X_2878_ _0630_ _0691_ u_bits.i_op1\[21\] _0692_ _0533_ _0658_ vssd1 vssd1 vccd1 vccd1
+ _0693_ sky130_fd_sc_hd__mux4_1
X_5597_ clknet_leaf_35_i_clk _0244_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[14\] sky130_fd_sc_hd__dfxtp_1
X_4548_ _1130_ _2006_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__nor2_1
X_4479_ u_muldiv.quotient_msk\[31\] _1210_ _1913_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__a21o_1
X_3850_ _0751_ _1345_ _0711_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__o21a_1
X_2801_ _0470_ _0615_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__xnor2_4
X_3781_ _0908_ _1503_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__nor2_1
X_5520_ clknet_leaf_13_i_clk _0168_ vssd1 vssd1 vccd1 vccd1 csr_data\[4\] sky130_fd_sc_hd__dfxtp_1
X_2732_ _0532_ _0544_ _0545_ _0546_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__o211a_1
X_5451_ clknet_leaf_9_i_clk _0099_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2663_ _0476_ _0477_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__nand2_1
X_5382_ clknet_leaf_48_i_clk _0030_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[14\] sky130_fd_sc_hd__dfxtp_2
X_4402_ u_bits.i_op2\[15\] _1906_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__or2_1
X_4333_ u_muldiv.divisor\[33\] _1838_ _1843_ u_muldiv.divisor\[34\] _1854_ vssd1 vssd1
+ vccd1 vccd1 _0199_ sky130_fd_sc_hd__a221o_1
X_4264_ _1806_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__clkbuf_1
X_3215_ _0962_ _0990_ _1013_ _0966_ _1014_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__o221a_1
X_4195_ u_wr_mux.i_reg_data2\[15\] i_reg_data2[15] _1767_ vssd1 vssd1 vccd1 vccd1
+ _1771_ sky130_fd_sc_hd__mux2_1
X_3146_ _0617_ _0639_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__and3_1
X_3077_ _0692_ u_bits.i_op2\[23\] _0634_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__a21o_1
X_5718_ clknet_leaf_24_i_clk _0361_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3979_ _0923_ _0831_ _1639_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__mux2_1
X_5649_ clknet_leaf_10_i_clk _0293_ vssd1 vssd1 vccd1 vccd1 op_cnt\[1\] sky130_fd_sc_hd__dfxtp_1
X_3000_ _0810_ _0811_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__and2_2
X_4951_ _1206_ _2309_ _2310_ _1828_ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__o31a_1
X_4882_ _2275_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__clkbuf_1
X_3902_ _1602_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__clkbuf_1
X_3833_ _1106_ csr_data\[17\] _1552_ _1124_ vssd1 vssd1 vccd1 vccd1 o_result[17] sky130_fd_sc_hd__o211a_2
X_3764_ _1487_ _0776_ _1267_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__a21oi_1
X_2715_ _0456_ _0529_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__xnor2_1
X_5503_ clknet_leaf_43_i_clk _0151_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_3695_ _1274_ _1422_ _1423_ _0624_ _1147_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__o32a_1
X_2646_ _0460_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__buf_2
X_5434_ clknet_leaf_1_i_clk _0082_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[25\] sky130_fd_sc_hd__dfxtp_4
X_5365_ clknet_leaf_39_i_clk _0013_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[61\] sky130_fd_sc_hd__dfxtp_1
X_5296_ u_muldiv.divisor\[10\] _2614_ _2615_ u_muldiv.divisor\[11\] vssd1 vssd1 vccd1
+ vccd1 _0401_ sky130_fd_sc_hd__a22o_1
X_4316_ u_muldiv.on_wait vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__clkinv_4
X_4247_ _1797_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
X_4178_ o_wdata[7] i_reg_data2[7] _1756_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__mux2_1
X_3129_ u_bits.i_op1\[25\] u_muldiv.add_prev\[25\] _0452_ vssd1 vssd1 vccd1 vccd1
+ _0935_ sky130_fd_sc_hd__mux2_2
X_3480_ o_wdata[6] u_wr_mux.i_reg_data2\[22\] _1224_ vssd1 vssd1 vccd1 vccd1 _1231_
+ sky130_fd_sc_hd__mux2_1
X_5150_ _0646_ _2362_ _2492_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__nand3_1
X_4101_ _1711_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__clkbuf_4
X_5081_ _2385_ _2428_ _0776_ vssd1 vssd1 vccd1 vccd1 _2430_ sky130_fd_sc_hd__a21o_1
X_4032_ u_bits.i_op2\[18\] u_bits.i_op2\[16\] _1657_ vssd1 vssd1 vccd1 vccd1 _1679_
+ sky130_fd_sc_hd__mux2_1
X_4934_ _2292_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__clkbuf_4
X_4865_ _2161_ _2261_ u_muldiv.o_div\[27\] vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__a21oi_1
X_4796_ _2167_ _2206_ u_muldiv.o_div\[13\] vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__a21oi_1
X_3816_ _0629_ _1530_ _0955_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__a21oi_1
X_3747_ _0670_ _0695_ _0642_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__a21oi_1
X_3678_ _1406_ _1258_ _0926_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__o22a_1
X_5417_ clknet_leaf_52_i_clk _0065_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[8\] sky130_fd_sc_hd__dfxtp_4
X_5348_ _1162_ _2628_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__nor2_1
X_5279_ _0699_ _2594_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__nor2_1
X_2980_ _0783_ _0792_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__or2b_1
X_4650_ u_muldiv.divisor\[7\] u_muldiv.dividend\[7\] vssd1 vssd1 vccd1 vccd1 _2073_
+ sky130_fd_sc_hd__and2b_1
X_3601_ _0730_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__clkbuf_2
X_4581_ _0993_ _2007_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__nor2_1
X_3532_ _0831_ _0917_ _0926_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__o22a_1
X_3463_ u_wr_mux.i_reg_data2\[14\] o_wdata[6] _0718_ vssd1 vssd1 vccd1 vccd1 _1222_
+ sky130_fd_sc_hd__mux2_1
X_5202_ _2120_ _2528_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__nor2_1
X_5133_ _2458_ _2093_ vssd1 vssd1 vccd1 vccd1 _2477_ sky130_fd_sc_hd__or2_1
X_3394_ _1104_ _1105_ _1167_ _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__o31a_1
X_5064_ u_muldiv.dividend\[12\] _2403_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__xor2_1
X_4015_ _1665_ _1666_ _1667_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__a21o_1
X_4917_ u_muldiv.quotient_msk\[25\] _2282_ _2283_ u_muldiv.quotient_msk\[26\] vssd1
+ vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__a22o_1
X_4848_ _2181_ _2246_ _2248_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__a21oi_1
X_4779_ u_muldiv.o_div\[9\] _2186_ u_muldiv.o_div\[10\] vssd1 vssd1 vccd1 vccd1 _2193_
+ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_2_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5751_ clknet_leaf_25_i_clk _0394_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2963_ u_bits.i_op1\[13\] vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__clkbuf_4
X_4702_ _2124_ u_muldiv.divisor\[26\] _2123_ u_muldiv.dividend\[27\] vssd1 vssd1 vccd1
+ vccd1 _2125_ sky130_fd_sc_hd__a2bb2o_1
X_5682_ clknet_leaf_32_i_clk _0325_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[28\] sky130_fd_sc_hd__dfxtp_1
X_2894_ _0708_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__inv_2
X_4633_ u_muldiv.divisor\[6\] u_muldiv.dividend\[6\] vssd1 vssd1 vccd1 vccd1 _2056_
+ sky130_fd_sc_hd__and2b_1
X_4564_ _2008_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__clkbuf_1
X_3515_ _0785_ _1250_ u_bits.i_op1\[10\] _1251_ _0778_ _0783_ vssd1 vssd1 vccd1 vccd1
+ _1252_ sky130_fd_sc_hd__mux4_1
X_4495_ u_muldiv.mul\[7\] u_muldiv.mul\[8\] _1978_ vssd1 vssd1 vccd1 vccd1 _1979_
+ sky130_fd_sc_hd__mux2_1
X_3446_ i_flush _1212_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__nor2_1
X_3377_ _1157_ vssd1 vssd1 vccd1 vccd1 o_add[12] sky130_fd_sc_hd__inv_2
X_5116_ _2459_ _2461_ _2288_ vssd1 vssd1 vccd1 vccd1 _2462_ sky130_fd_sc_hd__mux2_1
X_5047_ u_muldiv.on_wait _2397_ _2398_ vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__and3_1
X_3300_ _1073_ _1075_ _1076_ _1072_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__a31o_2
X_4280_ csr_data\[22\] i_csr_data[22] _1811_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__mux2_1
X_3231_ _1029_ u_bits.i_op1\[27\] _0689_ _0943_ _0778_ _0779_ vssd1 vssd1 vccd1 vccd1
+ _1030_ sky130_fd_sc_hd__mux4_1
X_3162_ _0934_ _0935_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__o21ai_2
X_3093_ _0895_ _0896_ _0900_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__a21o_1
X_5803_ clknet_leaf_34_i_clk _0445_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[51\] sky130_fd_sc_hd__dfxtp_1
X_3995_ _1406_ _1376_ _1639_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__mux2_1
X_5734_ clknet_leaf_18_i_clk _0377_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[18\]
+ sky130_fd_sc_hd__dfxtp_2
X_2946_ _0754_ _0757_ _0758_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__mux2_1
X_5665_ clknet_leaf_29_i_clk _0308_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[11\] sky130_fd_sc_hd__dfxtp_1
X_2877_ u_bits.i_op1\[23\] vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__clkbuf_4
X_4616_ u_muldiv.dividend\[15\] u_muldiv.divisor\[15\] vssd1 vssd1 vccd1 vccd1 _2039_
+ sky130_fd_sc_hd__and2b_1
X_5596_ clknet_leaf_36_i_clk _0243_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[13\] sky130_fd_sc_hd__dfxtp_1
X_4547_ _1214_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__buf_2
X_4478_ u_muldiv.divisor\[62\] _1210_ _1970_ u_bits.i_op2\[31\] vssd1 vssd1 vccd1
+ vccd1 _0228_ sky130_fd_sc_hd__a22o_1
X_3429_ op_cnt\[1\] _1197_ _1198_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_20_i_clk clknet_2_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2800_ _0496_ _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__nand2_2
X_3780_ _1110_ _1085_ _1500_ _1248_ _1502_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__a221o_1
X_2731_ _0530_ _0531_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_35_i_clk clknet_2_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5450_ clknet_leaf_9_i_clk _0098_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2662_ u_bits.i_op1\[18\] u_muldiv.add_prev\[18\] _0451_ vssd1 vssd1 vccd1 vccd1
+ _0477_ sky130_fd_sc_hd__mux2_1
X_4401_ u_muldiv.divisor\[46\] _1867_ _1887_ u_muldiv.divisor\[47\] _1909_ vssd1 vssd1
+ vccd1 vccd1 _0212_ sky130_fd_sc_hd__a221o_1
X_5381_ clknet_leaf_48_i_clk _0029_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[13\] sky130_fd_sc_hd__dfxtp_2
X_4332_ _1851_ _1853_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__nor2_1
X_4263_ csr_data\[14\] i_csr_data[14] _1800_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__mux2_1
X_3214_ _0987_ _0988_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__nand2_1
X_4194_ _1770_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__clkbuf_1
X_3145_ _0943_ u_bits.i_op2\[25\] vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__nand2_1
X_3076_ _0858_ _0865_ _0869_ _0884_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__or4_1
X_3978_ _1635_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__buf_2
X_2929_ _0633_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__buf_2
X_5717_ clknet_leaf_24_i_clk _0360_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_5648_ clknet_leaf_10_i_clk _0292_ vssd1 vssd1 vccd1 vccd1 op_cnt\[0\] sky130_fd_sc_hd__dfxtp_1
X_5579_ clknet_leaf_9_i_clk _0226_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_4950_ _2295_ _2308_ _1255_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__a21oi_1
X_4881_ u_muldiv.o_div\[30\] _2274_ _2244_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__mux2_1
X_3901_ _1310_ i_op1[4] _1599_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__mux2_1
X_3832_ _1541_ _1551_ _0446_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__a21o_1
X_5502_ clknet_leaf_43_i_clk _0150_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_3763_ u_bits.i_op2\[13\] vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__clkbuf_4
X_2714_ _0459_ u_bits.i_op2\[2\] u_bits.i_op1\[2\] _0463_ vssd1 vssd1 vccd1 vccd1
+ _0529_ sky130_fd_sc_hd__a22o_1
X_3694_ u_bits.i_op2\[8\] _0785_ _1272_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__a21oi_1
X_2645_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__buf_2
X_5433_ clknet_leaf_0_i_clk _0081_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[24\] sky130_fd_sc_hd__dfxtp_2
X_5364_ clknet_leaf_34_i_clk _0012_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[60\] sky130_fd_sc_hd__dfxtp_1
X_4315_ _1835_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__buf_2
X_5295_ u_muldiv.divisor\[9\] _2614_ _2615_ u_muldiv.divisor\[10\] vssd1 vssd1 vccd1
+ vccd1 _0400_ sky130_fd_sc_hd__a22o_1
X_4246_ csr_data\[6\] i_csr_data[6] _1789_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__mux2_1
X_4177_ _1761_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__clkbuf_1
X_3128_ _0458_ _0933_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__xnor2_4
X_3059_ _0692_ u_bits.i_op2\[23\] _0867_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__a21oi_1
X_5080_ _0776_ _2293_ _2428_ vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__nand3_1
X_4100_ _1722_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__clkbuf_1
X_4031_ _1665_ _1677_ _1678_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__a21o_1
X_4933_ _0917_ _0791_ _2293_ u_muldiv.on_wait vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__a31o_1
X_4864_ u_muldiv.quotient_msk\[27\] _2258_ _2229_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__mux2_1
X_4795_ u_muldiv.quotient_msk\[13\] _2201_ _2156_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__mux2_1
X_3815_ _0628_ _1529_ _1532_ _1535_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__or4_1
X_3746_ _0788_ _1470_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__or2_1
X_5416_ clknet_leaf_46_i_clk _0064_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[7\] sky130_fd_sc_hd__dfxtp_1
X_3677_ _1406_ _1258_ _0867_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__a21oi_1
X_5347_ _1163_ _2628_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__nor2_1
X_5278_ _2607_ _2608_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__xnor2_1
X_4229_ _1788_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_1
X_3600_ _1106_ csr_data\[2\] _1124_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__o21ai_1
X_4580_ _2014_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__clkbuf_1
X_3531_ _0831_ _0917_ _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__a21oi_1
X_3462_ _1221_ vssd1 vssd1 vccd1 vccd1 o_wdata[13] sky130_fd_sc_hd__buf_2
X_5201_ _0904_ _2293_ _2537_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__and3_1
X_3393_ _1095_ _1099_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__nand2_1
X_5132_ u_muldiv.dividend\[18\] _2468_ vssd1 vssd1 vccd1 vccd1 _2476_ sky130_fd_sc_hd__xor2_1
X_5063_ _2413_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__clkbuf_1
X_4014_ u_bits.i_op2\[11\] _1663_ _1651_ i_op2[11] vssd1 vssd1 vccd1 vccd1 _1667_
+ sky130_fd_sc_hd__a22o_1
X_4916_ u_muldiv.quotient_msk\[24\] _2282_ _2283_ u_muldiv.quotient_msk\[25\] vssd1
+ vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__a22o_1
X_4847_ _2161_ _2247_ u_muldiv.o_div\[23\] vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__a21oi_1
X_4778_ _2181_ _2190_ _2192_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__a21oi_1
X_3729_ _1333_ csr_data\[10\] _1388_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__o21ai_1
X_5750_ clknet_leaf_24_i_clk _0393_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2962_ _0772_ _0773_ _0774_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__mux2_2
X_5681_ clknet_leaf_31_i_clk _0324_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[27\] sky130_fd_sc_hd__dfxtp_1
X_4701_ _2123_ u_muldiv.dividend\[27\] u_muldiv.dividend\[26\] vssd1 vssd1 vccd1 vccd1
+ _2124_ sky130_fd_sc_hd__o21ai_1
X_4632_ u_muldiv.dividend\[7\] u_muldiv.divisor\[7\] vssd1 vssd1 vccd1 vccd1 _2055_
+ sky130_fd_sc_hd__and2b_1
X_2893_ _0695_ _0706_ _0707_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__mux2_1
X_4563_ o_add[16] _2004_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__and2_1
X_4494_ _1583_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__clkbuf_4
X_3514_ u_bits.i_op1\[11\] vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__buf_4
X_3445_ _1204_ i_alu_ctrl[1] _1202_ _1211_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__o2bb2a_1
X_3376_ _1153_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__nand2_4
X_5115_ _0653_ _2460_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__xnor2_1
X_5046_ _2051_ _2077_ _2050_ vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__o21ai_1
X_3230_ u_bits.i_op1\[28\] vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__clkbuf_4
X_3161_ _0898_ _0899_ _0934_ _0935_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__a22o_1
X_3092_ _0898_ _0899_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__xnor2_1
X_5802_ clknet_leaf_39_i_clk _0444_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[50\] sky130_fd_sc_hd__dfxtp_1
X_3994_ _1641_ _1650_ _1652_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__a21o_1
X_5733_ clknet_leaf_18_i_clk _0376_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[17\]
+ sky130_fd_sc_hd__dfxtp_2
X_2945_ u_bits.i_op2\[2\] vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__clkbuf_4
X_5664_ clknet_leaf_28_i_clk _0307_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[10\] sky130_fd_sc_hd__dfxtp_1
X_2876_ u_bits.i_op1\[22\] vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__buf_4
X_4615_ u_muldiv.divisor\[18\] _2037_ u_muldiv.dividend\[18\] vssd1 vssd1 vccd1 vccd1
+ _2038_ sky130_fd_sc_hd__or3b_1
X_5595_ clknet_leaf_36_i_clk _0242_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[12\] sky130_fd_sc_hd__dfxtp_1
X_4546_ _2005_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
X_4477_ _1868_ _1969_ _1833_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__a21oi_1
X_3428_ u_muldiv.i_is_div vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__buf_6
X_3359_ _0594_ _1144_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__xor2_4
X_5029_ _2052_ _2371_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__nand2_1
Xclkbuf_2_1__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_1_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2730_ _0526_ _0527_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__nand2_1
X_2661_ _0457_ _0475_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__xnor2_1
X_4400_ _1907_ _1908_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__nor2_1
X_5380_ clknet_leaf_48_i_clk _0028_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[12\] sky130_fd_sc_hd__dfxtp_2
X_4331_ _0923_ _0915_ _1852_ _1832_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__a31o_1
X_4262_ _1805_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__clkbuf_1
X_3213_ _0964_ _0991_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__nand2_1
X_4193_ u_wr_mux.i_reg_data2\[14\] i_reg_data2[14] _1767_ vssd1 vssd1 vccd1 vccd1
+ _1770_ sky130_fd_sc_hd__mux2_1
X_3144_ _0947_ _0948_ _0707_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__mux2_1
X_3075_ _0643_ _0878_ _0883_ _0800_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__o211a_1
X_3977_ _0831_ _1637_ _1638_ i_op2[0] _1640_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__a221o_1
X_5716_ clknet_leaf_36_i_clk _0359_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_2928_ _0719_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__buf_2
X_5647_ clknet_leaf_8_i_clk _0000_ vssd1 vssd1 vccd1 vccd1 u_muldiv.i_on_end sky130_fd_sc_hd__dfxtp_2
X_2859_ _0673_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__clkbuf_4
X_5578_ clknet_leaf_9_i_clk _0225_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_4529_ _1996_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__clkbuf_1
X_4880_ _2271_ _2272_ _2273_ _1841_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__a22o_1
X_3900_ _1601_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__clkbuf_1
X_3831_ _0749_ o_add[17] _1549_ _1550_ _0453_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__a221o_1
X_3762_ _0759_ _1485_ _0824_ _0765_ _0920_ _0643_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__mux4_1
X_5501_ clknet_leaf_43_i_clk _0149_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_2713_ _0526_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__nor2_1
X_3693_ _0908_ _1421_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__nor2_1
X_2644_ u_mux.i_group_mux vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__inv_2
X_5432_ clknet_leaf_0_i_clk _0080_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[23\] sky130_fd_sc_hd__dfxtp_4
X_5363_ clknet_leaf_39_i_clk _0011_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[59\] sky130_fd_sc_hd__dfxtp_1
X_4314_ u_muldiv.divisor\[32\] _1829_ _1833_ _0831_ _1837_ vssd1 vssd1 vccd1 vccd1
+ _0197_ sky130_fd_sc_hd__o221a_1
X_5294_ _1842_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__buf_2
X_4245_ _1796_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
X_4176_ o_wdata[6] i_reg_data2[6] _1756_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__mux2_1
X_3127_ _0461_ u_bits.i_op2\[25\] _0465_ u_bits.i_op1\[25\] vssd1 vssd1 vccd1 vccd1
+ _0933_ sky130_fd_sc_hd__a22o_1
X_3058_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_34_i_clk clknet_2_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_49_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4030_ u_bits.i_op2\[16\] _1663_ _1675_ i_op2[16] vssd1 vssd1 vccd1 vccd1 _1678_
+ sky130_fd_sc_hd__a22o_1
X_4932_ _2292_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__buf_2
X_4863_ u_muldiv.o_div\[27\] _2170_ _2258_ _2196_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__a31o_1
X_4794_ _2170_ u_muldiv.o_div\[13\] _2201_ _2196_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__a31o_1
X_3814_ _0672_ _1533_ _1534_ _0800_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__o211a_1
X_3745_ _1253_ _1261_ _0668_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__mux2_1
X_3676_ u_bits.i_op2\[7\] vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__buf_4
X_5415_ clknet_leaf_49_i_clk _0063_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[6\] sky130_fd_sc_hd__dfxtp_4
X_5346_ _1155_ _2628_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__nor2_1
X_5277_ _2137_ _2144_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__nor2_1
X_4228_ u_wr_mux.i_reg_data2\[31\] i_reg_data2[31] _1778_ vssd1 vssd1 vccd1 vccd1
+ _1788_ sky130_fd_sc_hd__mux2_1
X_4159_ u_bits.i_sra i_alu_ctrl[3] _1745_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__mux2_1
X_3530_ _0867_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__clkbuf_4
X_3461_ u_wr_mux.i_reg_data2\[13\] o_wdata[5] _0718_ vssd1 vssd1 vccd1 vccd1 _1221_
+ sky130_fd_sc_hd__mux2_1
X_5200_ _2295_ _2537_ _0904_ vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__a21oi_1
X_3392_ _1095_ _1099_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__nor2_1
X_5131_ _2475_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__clkbuf_1
X_5062_ u_muldiv.dividend\[11\] _2412_ _2378_ vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__mux2_1
X_4013_ u_bits.i_op2\[12\] _1445_ _1657_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__mux2_1
X_4915_ u_muldiv.quotient_msk\[23\] _2282_ _2283_ u_muldiv.quotient_msk\[24\] vssd1
+ vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__a22o_1
X_4846_ u_muldiv.quotient_msk\[23\] _2241_ _2229_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__mux2_1
X_4777_ _2167_ _2191_ u_muldiv.o_div\[9\] vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__a21oi_1
X_3728_ _1331_ _1451_ _1453_ _1454_ _1357_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__o221a_1
X_3659_ _1309_ _1314_ _1312_ _1306_ _0669_ _0920_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__mux4_1
X_5329_ _2625_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__clkbuf_1
X_2961_ _0659_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__clkbuf_4
X_5680_ clknet_leaf_31_i_clk _0323_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[26\] sky130_fd_sc_hd__dfxtp_1
X_4700_ u_muldiv.divisor\[27\] vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__inv_2
X_4631_ _2052_ _2053_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__nand2_1
X_2892_ _0524_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__clkbuf_4
X_4562_ _1162_ _2007_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__nor2_1
X_4493_ _1977_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_1
X_3513_ u_bits.i_op1\[9\] vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__buf_4
X_3444_ u_muldiv.i_on_wait vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__clkinv_2
X_3375_ _0578_ _1152_ _0607_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__nand3_1
X_5114_ _0654_ _2450_ _2385_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__o21ai_1
X_5045_ _2050_ _2051_ _2077_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__or3_1
X_4829_ u_muldiv.o_div\[20\] u_muldiv.o_div\[19\] _2226_ vssd1 vssd1 vccd1 vccd1 _2233_
+ sky130_fd_sc_hd__or3_2
X_3160_ _0962_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__and2_2
X_3091_ u_bits.i_op1\[24\] u_muldiv.add_prev\[24\] _0452_ vssd1 vssd1 vccd1 vccd1
+ _0899_ sky130_fd_sc_hd__mux2_1
X_5801_ clknet_leaf_35_i_clk _0443_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[49\] sky130_fd_sc_hd__dfxtp_1
X_5732_ clknet_leaf_18_i_clk _0375_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_3993_ _1376_ _1637_ _1651_ i_op2[5] vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__a22o_1
X_2944_ _0755_ _0756_ _0648_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__mux2_1
X_5663_ clknet_leaf_27_i_clk _0306_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[9\] sky130_fd_sc_hd__dfxtp_1
X_2875_ u_bits.i_op1\[24\] u_bits.i_op1\[25\] _0689_ u_bits.i_op1\[27\] _0650_ _0659_
+ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__mux4_1
X_4614_ u_muldiv.dividend\[19\] u_muldiv.divisor\[19\] vssd1 vssd1 vccd1 vccd1 _2037_
+ sky130_fd_sc_hd__and2b_1
X_5594_ clknet_leaf_36_i_clk _0241_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[11\] sky130_fd_sc_hd__dfxtp_1
X_4545_ o_add[1] _2004_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__and2_1
X_4476_ u_bits.i_op2\[29\] u_bits.i_op2\[30\] _1962_ vssd1 vssd1 vccd1 vccd1 _1969_
+ sky130_fd_sc_hd__or3_1
X_3427_ op_cnt\[2\] op_cnt\[3\] op_cnt\[4\] op_cnt\[5\] vssd1 vssd1 vccd1 vccd1 _1197_
+ sky130_fd_sc_hd__or4b_1
X_3358_ _0596_ _0597_ _1143_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__a21bo_1
X_3289_ _0832_ _0833_ _1083_ _0976_ _0825_ _0920_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__mux4_1
X_5028_ u_muldiv.dividend\[8\] _2361_ u_muldiv.dividend\[9\] vssd1 vssd1 vccd1 vccd1
+ _2381_ sky130_fd_sc_hd__o21ai_1
X_2660_ _0460_ u_bits.i_op2\[18\] u_bits.i_op1\[18\] _0464_ vssd1 vssd1 vccd1 vccd1
+ _0475_ sky130_fd_sc_hd__a22o_1
X_4330_ _1845_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__buf_2
X_4261_ csr_data\[13\] i_csr_data[13] _1800_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__mux2_1
X_3212_ _0739_ csr_data\[27\] _1012_ _0732_ vssd1 vssd1 vccd1 vccd1 o_result[27] sky130_fd_sc_hd__o211a_2
X_4192_ _1769_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__clkbuf_1
X_3143_ _0669_ _0793_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__nor2_1
X_3074_ _0879_ _0882_ _0642_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__a21bo_1
X_3976_ _1639_ _1635_ _1112_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__and3b_1
X_5715_ clknet_leaf_32_i_clk _0358_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_2927_ _0622_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__buf_2
X_5646_ clknet_leaf_11_i_clk _0002_ vssd1 vssd1 vccd1 vccd1 u_muldiv.i_on_wait sky130_fd_sc_hd__dfxtp_2
X_2858_ _0524_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__inv_2
X_5577_ clknet_leaf_9_i_clk _0224_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_2789_ _0592_ _0593_ _0596_ _0597_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__a22o_1
X_4528_ u_muldiv.mul\[23\] u_muldiv.mul\[24\] _1989_ vssd1 vssd1 vccd1 vccd1 _1996_
+ sky130_fd_sc_hd__mux2_1
X_4459_ u_bits.i_op2\[27\] _1955_ _1832_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__a21oi_1
X_3830_ _0629_ _1543_ _0955_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__a21oi_1
X_3761_ _1282_ _1288_ _0758_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__mux2_1
X_2712_ u_bits.i_op1\[3\] u_muldiv.add_prev\[3\] _0450_ vssd1 vssd1 vccd1 vccd1 _0527_
+ sky130_fd_sc_hd__mux2_1
X_5500_ clknet_leaf_43_i_clk _0148_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_3692_ _1110_ _0921_ _1418_ _1249_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__a221o_1
X_2643_ _0457_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__buf_6
X_5431_ clknet_leaf_0_i_clk _0079_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[22\] sky130_fd_sc_hd__dfxtp_4
X_5362_ clknet_leaf_40_i_clk _0010_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[58\] sky130_fd_sc_hd__dfxtp_1
X_4313_ _1834_ _1836_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__nand2_1
X_5293_ u_muldiv.divisor\[8\] _2614_ _2285_ u_muldiv.divisor\[9\] vssd1 vssd1 vccd1
+ vccd1 _0399_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_0_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4244_ csr_data\[5\] i_csr_data[5] _1789_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__mux2_1
X_4175_ _1760_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__clkbuf_1
X_3126_ _0739_ csr_data\[24\] _0932_ _0732_ vssd1 vssd1 vccd1 vccd1 o_result[24] sky130_fd_sc_hd__o211a_2
X_3057_ o_funct3[2] _0638_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__nand2_1
X_3959_ _1596_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__clkbuf_4
X_5629_ clknet_leaf_44_i_clk _0276_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_4931_ _2291_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__buf_2
X_4862_ u_muldiv.o_div\[26\] _2171_ _2259_ _2164_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__a22o_1
X_3813_ _0672_ _1266_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__nand2_1
X_4793_ _2204_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__clkbuf_1
X_3744_ _1468_ _1469_ _1336_ u_pc_sel.i_pc_next\[11\] vssd1 vssd1 vccd1 vccd1 o_result[11]
+ sky130_fd_sc_hd__a2bb2o_2
X_3675_ _1404_ _0864_ _0751_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__mux2_1
X_5414_ clknet_leaf_49_i_clk _0062_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[5\] sky130_fd_sc_hd__dfxtp_1
X_5345_ _1157_ _2628_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__nor2_1
X_5276_ _2136_ u_muldiv.dividend\[30\] _2135_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__a21oi_1
X_4227_ _1787_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__clkbuf_1
X_4158_ _1751_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__clkbuf_1
X_3109_ u_bits.i_op2\[2\] _0915_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__or2_2
X_4089_ u_pc_sel.i_pc_next\[5\] i_pc_next[5] _1712_ vssd1 vssd1 vccd1 vccd1 _1717_
+ sky130_fd_sc_hd__mux2_1
X_3460_ _1220_ vssd1 vssd1 vccd1 vccd1 o_wdata[12] sky130_fd_sc_hd__buf_2
X_3391_ _0616_ vssd1 vssd1 vccd1 vccd1 o_add[20] sky130_fd_sc_hd__inv_2
X_5130_ u_muldiv.dividend\[17\] _2474_ _2378_ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__mux2_1
X_5061_ _1208_ _2403_ _2404_ _2408_ _2411_ vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__a32o_1
X_4012_ _1635_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__buf_2
X_4914_ u_muldiv.quotient_msk\[22\] _2282_ _2283_ u_muldiv.quotient_msk\[23\] vssd1
+ vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__a22o_1
X_4845_ u_muldiv.o_div\[23\] _2170_ _2241_ _2196_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__a31o_1
X_4776_ u_muldiv.quotient_msk\[9\] _2186_ _2156_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__mux2_1
X_3727_ u_muldiv.mul\[10\] _1330_ _1400_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_33_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3658_ _1387_ _1389_ _1336_ u_pc_sel.i_pc_next\[5\] vssd1 vssd1 vccd1 vccd1 o_result[5]
+ sky130_fd_sc_hd__a2bb2o_2
X_3589_ _1274_ _1322_ _1323_ _0624_ _1130_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__o32a_1
X_5328_ u_muldiv.dividend\[0\] _2624_ _2152_ vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_48_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5259_ _1208_ _2583_ _2584_ _2591_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__a31o_1
X_2960_ u_bits.i_op1\[19\] _0645_ _0656_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__mux2_1
X_2891_ _0705_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__clkinv_2
X_4630_ u_muldiv.dividend\[8\] u_muldiv.divisor\[8\] vssd1 vssd1 vccd1 vccd1 _2053_
+ sky130_fd_sc_hd__or2b_1
X_4561_ _1163_ _2007_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__nor2_1
X_4492_ u_muldiv.mul\[6\] u_muldiv.mul\[7\] _1584_ vssd1 vssd1 vccd1 vccd1 _1977_
+ sky130_fd_sc_hd__mux2_1
X_3512_ _1248_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__clkbuf_4
X_3443_ _1204_ _1205_ _1210_ i_flush vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a211o_1
X_5113_ _2458_ _2089_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__xor2_1
X_3374_ _1155_ vssd1 vssd1 vccd1 vccd1 o_add[13] sky130_fd_sc_hd__inv_2
X_5044_ _2295_ _2394_ _1305_ vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__a21o_1
X_4828_ u_muldiv.o_div\[19\] _2226_ u_muldiv.o_div\[20\] vssd1 vssd1 vccd1 vccd1 _2232_
+ sky130_fd_sc_hd__o21ai_1
X_4759_ _2164_ _2175_ _2177_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__a21oi_1
X_3090_ _0458_ _0897_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__xnor2_2
X_3992_ _1595_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__buf_2
X_5800_ clknet_leaf_39_i_clk _0442_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[48\] sky130_fd_sc_hd__dfxtp_1
X_5731_ clknet_leaf_21_i_clk _0374_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_2943_ u_bits.i_op1\[27\] u_bits.i_op1\[28\] _0649_ vssd1 vssd1 vccd1 vccd1 _0756_
+ sky130_fd_sc_hd__mux2_1
X_5662_ clknet_leaf_26_i_clk _0305_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[8\] sky130_fd_sc_hd__dfxtp_1
X_2874_ u_bits.i_op1\[26\] vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__buf_4
X_4613_ u_muldiv.divisor\[19\] u_muldiv.dividend\[19\] vssd1 vssd1 vccd1 vccd1 _2036_
+ sky130_fd_sc_hd__or2b_1
X_5593_ clknet_leaf_36_i_clk _0240_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[10\] sky130_fd_sc_hd__dfxtp_1
X_4544_ _1583_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__clkbuf_4
X_4475_ u_muldiv.divisor\[61\] _1836_ _1946_ u_muldiv.divisor\[62\] _1968_ vssd1 vssd1
+ vccd1 vccd1 _0227_ sky130_fd_sc_hd__a221o_1
X_3426_ u_pc_sel.i_inst_branch _1191_ _1196_ u_pc_sel.i_inst_jal_jalr vssd1 vssd1
+ vccd1 vccd1 o_pc_select sky130_fd_sc_hd__a31o_2
X_3357_ _0568_ _0576_ _0598_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__a21o_1
X_5027_ u_muldiv.dividend\[9\] u_muldiv.dividend\[8\] _2361_ vssd1 vssd1 vccd1 vccd1
+ _2380_ sky130_fd_sc_hd__or3_1
X_3288_ _0699_ _0697_ _1029_ _0996_ _0651_ _0774_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__mux4_1
X_4260_ _1804_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_1
X_3211_ _0995_ _1011_ _0447_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__a21o_1
X_4191_ u_wr_mux.i_reg_data2\[13\] i_reg_data2[13] _1767_ vssd1 vssd1 vccd1 vccd1
+ _1769_ sky130_fd_sc_hd__mux2_1
X_3142_ _0787_ _0795_ _0758_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__mux2_1
X_3073_ _0880_ _0881_ _0696_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__mux2_1
X_3975_ _1198_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__clkbuf_4
X_5714_ clknet_leaf_33_i_clk _0357_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_2926_ _0728_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__buf_2
X_5645_ clknet_leaf_9_i_clk _0001_ vssd1 vssd1 vccd1 vccd1 o_ready sky130_fd_sc_hd__dfxtp_2
X_2857_ _0642_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__buf_2
X_5576_ clknet_leaf_9_i_clk _0223_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_2788_ _0587_ _0588_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__nand2_1
X_4527_ _1995_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__clkbuf_1
X_4458_ u_bits.i_op2\[26\] _1942_ _1951_ _1845_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__o31a_1
X_3409_ _1135_ _1142_ _1147_ _1179_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__and4_1
X_4389_ _1868_ _1899_ _1487_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__a21oi_1
X_3760_ _1483_ _1484_ _0730_ u_pc_sel.i_pc_next\[12\] vssd1 vssd1 vccd1 vccd1 o_result[12]
+ sky130_fd_sc_hd__a2bb2o_2
X_2711_ _0457_ _0525_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__xnor2_1
X_5430_ clknet_leaf_1_i_clk _0078_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[21\] sky130_fd_sc_hd__dfxtp_4
X_3691_ u_bits.i_op2\[8\] _0785_ _0637_ _1419_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__o22a_1
X_2642_ _0456_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__buf_6
X_5361_ clknet_leaf_39_i_clk _0009_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[57\] sky130_fd_sc_hd__dfxtp_1
X_5292_ u_muldiv.divisor\[7\] _2614_ _2285_ u_muldiv.divisor\[8\] vssd1 vssd1 vccd1
+ vccd1 _0398_ sky130_fd_sc_hd__a22o_1
X_4312_ _1835_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__buf_2
X_4243_ _1795_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
X_4174_ o_wdata[5] i_reg_data2[5] _1756_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__mux2_1
X_3125_ _0892_ _0931_ _0447_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__a21o_1
X_3056_ _0643_ _0864_ _0711_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__o21a_1
X_3958_ _1631_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__clkbuf_1
X_3889_ i_flush i_reset_n o_ready vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__and3b_1
X_2909_ _0461_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__clkbuf_4
X_5628_ clknet_leaf_44_i_clk _0275_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_5559_ clknet_leaf_7_i_clk _0206_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_4930_ _0620_ _0702_ vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__and2b_1
X_4861_ _2165_ _2257_ _2258_ _1842_ u_muldiv.quotient_msk\[26\] vssd1 vssd1 vccd1
+ vccd1 _2259_ sky130_fd_sc_hd__a32o_1
X_3812_ _0660_ _0664_ _0667_ _0678_ _0825_ _0707_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__mux4_1
X_4792_ u_muldiv.o_div\[12\] _2203_ _2154_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__mux2_1
X_3743_ _1333_ csr_data\[11\] _1388_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__o21ai_1
X_3674_ _1339_ _1343_ _1341_ _1337_ _0669_ _0920_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__mux4_1
X_5413_ clknet_leaf_49_i_clk _0061_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[4\] sky130_fd_sc_hd__dfxtp_2
X_5344_ _1150_ _2628_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__nor2_1
X_5275_ u_muldiv.dividend\[31\] _2601_ _2605_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__a21o_1
X_4226_ u_wr_mux.i_reg_data2\[30\] i_reg_data2[30] _1778_ vssd1 vssd1 vccd1 vccd1
+ _1787_ sky130_fd_sc_hd__mux2_1
X_4157_ alu_ctrl\[2\] i_alu_ctrl[2] _1745_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__mux2_1
X_3108_ u_bits.i_op2\[0\] u_bits.i_op2\[1\] vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__or2_1
X_4088_ _1716_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__clkbuf_1
X_3039_ _0458_ _0848_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__xnor2_1
X_3390_ _0483_ _1165_ vssd1 vssd1 vccd1 vccd1 o_add[18] sky130_fd_sc_hd__xnor2_4
X_5060_ _2375_ _2410_ _1207_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__a21oi_1
X_4011_ _1641_ _1662_ _1664_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__a21o_1
X_4913_ u_muldiv.quotient_msk\[21\] _2282_ _2283_ u_muldiv.quotient_msk\[22\] vssd1
+ vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__a22o_1
X_4844_ _2245_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__clkbuf_1
X_4775_ _2165_ u_muldiv.o_div\[9\] _2186_ _1913_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__a31o_1
X_3726_ u_muldiv.mul\[42\] _1325_ _1452_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__a21oi_1
X_3657_ _1106_ csr_data\[5\] _1388_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__o21ai_1
X_3588_ _0923_ _1255_ _1272_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__a21oi_1
X_5327_ _0917_ _1880_ _2623_ _1841_ vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__a22o_1
X_5258_ _2586_ _2587_ _2590_ _1827_ vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__o211a_1
X_5189_ _2031_ _2105_ _2106_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__nor3_1
X_4209_ _1711_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__clkbuf_4
X_2890_ _0696_ _0701_ _0704_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__o21a_1
X_4560_ _1155_ _2007_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__nor2_1
X_4491_ _1976_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__clkbuf_1
X_3511_ _0710_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__clkinv_2
X_3442_ _1209_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__buf_4
X_3373_ _0577_ _1154_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__xor2_4
X_5112_ _2039_ _2083_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__or2_1
X_5043_ _1305_ _2362_ _2394_ vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__nand3_1
X_4827_ _2181_ _2228_ _2231_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__a21oi_1
X_4758_ _2167_ _2176_ u_muldiv.o_div\[5\] vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__a21oi_1
X_4689_ _2109_ _2111_ vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__nand2_1
X_3709_ _0714_ _1435_ _1436_ _0624_ _1145_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_32_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3991_ u_bits.i_op2\[6\] _0688_ _1639_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__mux2_1
X_5730_ clknet_leaf_20_i_clk _0373_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_2942_ u_bits.i_op1\[25\] _0689_ _0649_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__mux2_1
X_5661_ clknet_leaf_27_i_clk _0304_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[7\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_47_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2873_ _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__buf_4
X_4612_ _2032_ _2033_ _2034_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__a21o_1
X_5592_ clknet_leaf_36_i_clk _0239_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[9\] sky130_fd_sc_hd__dfxtp_1
X_4543_ _2003_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
X_4474_ _1832_ _1967_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__nor2_1
X_3425_ _1192_ _1195_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__nand2_1
X_3356_ _1142_ vssd1 vssd1 vccd1 vccd1 o_add[6] sky130_fd_sc_hd__inv_2
X_3287_ _0644_ _1081_ _0712_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__o21a_1
X_5026_ _2379_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__clkbuf_1
X_4190_ _1768_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__clkbuf_1
X_3210_ _0750_ o_add[27] _0997_ _1010_ _0804_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__a221o_1
X_3141_ _0784_ _0780_ _0945_ _0775_ _0825_ _0920_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__mux4_2
X_3072_ u_bits.i_op1\[3\] u_bits.i_op1\[2\] _0791_ u_bits.i_op1\[0\] _0657_ _0648_
+ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__mux4_1
X_3974_ _1595_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__clkbuf_4
X_5713_ clknet_leaf_32_i_clk _0356_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_2925_ _0736_ _0738_ vssd1 vssd1 vccd1 vccd1 o_add[21] sky130_fd_sc_hd__xnor2_4
X_2856_ _0652_ _0660_ _0664_ _0667_ _0669_ _0670_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__mux4_2
X_5644_ clknet_leaf_39_i_clk _0291_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_5575_ clknet_leaf_9_i_clk _0222_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_2787_ _0582_ _0583_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__nor2_1
X_4526_ u_muldiv.mul\[22\] u_muldiv.mul\[23\] _1989_ vssd1 vssd1 vccd1 vccd1 _1995_
+ sky130_fd_sc_hd__mux2_1
X_4457_ u_muldiv.divisor\[57\] _1836_ _1946_ u_muldiv.divisor\[58\] _1954_ vssd1 vssd1
+ vccd1 vccd1 _0223_ sky130_fd_sc_hd__a221o_1
X_3408_ _1128_ _1130_ _1137_ _1178_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__and4_1
X_4388_ u_bits.i_op2\[12\] _1895_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__or2_1
X_3339_ _1125_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__nand2_4
X_5009_ _1258_ _2362_ _2363_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__nand3_1
X_2710_ _0460_ _0524_ u_bits.i_op1\[3\] _0464_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__a22o_1
X_3690_ u_bits.i_op2\[8\] _0785_ _1267_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__a21oi_1
X_2641_ _0455_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__clkbuf_16
X_5360_ clknet_leaf_39_i_clk _0008_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[56\] sky130_fd_sc_hd__dfxtp_1
X_5291_ u_muldiv.divisor\[6\] _2614_ _2285_ u_muldiv.divisor\[7\] vssd1 vssd1 vccd1
+ vccd1 _0397_ sky130_fd_sc_hd__a22o_1
X_4311_ _1207_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__buf_4
X_4242_ csr_data\[4\] i_csr_data[4] _1789_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__mux2_1
X_4173_ _1759_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__clkbuf_1
X_3124_ _0750_ o_add[24] _0907_ _0930_ _0804_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__a221o_1
X_3055_ _0860_ _0863_ _0673_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__mux2_1
X_3957_ _0702_ i_op1[31] _1621_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__mux2_1
X_2908_ _0722_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__buf_2
X_3888_ _1593_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__clkbuf_1
X_5627_ clknet_leaf_44_i_clk _0274_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_2839_ u_bits.i_op1\[15\] vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__buf_4
X_5558_ clknet_leaf_7_i_clk _0205_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_4509_ u_muldiv.mul\[14\] u_muldiv.mul\[15\] _1978_ vssd1 vssd1 vccd1 vccd1 _1986_
+ sky130_fd_sc_hd__mux2_1
X_5489_ clknet_leaf_51_i_clk _0137_ vssd1 vssd1 vccd1 vccd1 o_wdata[7] sky130_fd_sc_hd__dfxtp_4
X_4860_ u_muldiv.o_div\[25\] u_muldiv.o_div\[26\] _2250_ vssd1 vssd1 vccd1 vccd1 _2258_
+ sky130_fd_sc_hd__or3_1
X_3811_ u_bits.i_op2\[16\] _0653_ _0637_ _1531_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__o22a_1
X_4791_ _1835_ _2200_ _2201_ _2202_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__a31o_1
X_3742_ _1331_ _1464_ _1466_ _1467_ _1357_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__o221a_1
X_3673_ _1402_ _1403_ _1336_ u_pc_sel.i_pc_next\[6\] vssd1 vssd1 vccd1 vccd1 o_result[6]
+ sky130_fd_sc_hd__a2bb2o_2
X_5412_ clknet_leaf_4_i_clk _0060_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[3\] sky130_fd_sc_hd__dfxtp_1
X_5343_ _1151_ _2628_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__nor2_1
X_5274_ u_muldiv.dividend\[31\] _2601_ _1835_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__o21ai_1
X_4225_ _1786_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__clkbuf_1
X_4156_ _1750_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__clkbuf_1
X_3107_ _0642_ _0625_ _0799_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__and3_2
X_4087_ u_pc_sel.i_pc_next\[4\] i_pc_next[4] _1712_ vssd1 vssd1 vccd1 vccd1 _1716_
+ sky130_fd_sc_hd__mux2_1
X_3038_ _0461_ u_bits.i_op2\[23\] _0465_ u_bits.i_op1\[23\] vssd1 vssd1 vccd1 vccd1
+ _0848_ sky130_fd_sc_hd__a22o_1
X_4989_ u_muldiv.dividend\[6\] _2336_ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__or2_1
X_4010_ _1445_ _1663_ _1651_ i_op2[10] vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__a22o_1
X_4912_ u_muldiv.quotient_msk\[20\] _2282_ _2283_ u_muldiv.quotient_msk\[21\] vssd1
+ vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__a22o_1
X_4843_ u_muldiv.o_div\[22\] _2243_ _2244_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__mux2_1
X_4774_ _2189_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__clkbuf_1
X_3725_ u_muldiv.dividend\[10\] _1326_ _1327_ u_muldiv.o_div\[10\] _1383_ vssd1 vssd1
+ vccd1 vccd1 _1452_ sky130_fd_sc_hd__a221o_1
X_3656_ _0731_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__clkbuf_2
X_3587_ _1249_ _1317_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__a21oi_1
X_5326_ _2063_ _2622_ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__nand2_1
X_5257_ _2288_ _2589_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__nand2_1
X_4208_ _1777_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__clkbuf_1
X_5188_ _2031_ _2105_ _2106_ _2120_ vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__o22a_1
X_4139_ _1741_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__clkbuf_1
X_3510_ _0620_ _1170_ _1246_ _0625_ _0619_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__o2111ai_2
X_4490_ u_muldiv.mul\[5\] u_muldiv.mul\[6\] _1584_ vssd1 vssd1 vccd1 vccd1 _1976_
+ sky130_fd_sc_hd__mux2_1
X_3441_ _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__buf_4
X_3372_ _0519_ _1153_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__nand2_1
X_5111_ u_muldiv.dividend\[16\] _2444_ vssd1 vssd1 vccd1 vccd1 _2457_ sky130_fd_sc_hd__xor2_1
X_5042_ u_bits.i_op1\[9\] _2386_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__or2_2
X_4826_ _2161_ _2230_ u_muldiv.o_div\[19\] vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__a21oi_1
X_4757_ u_muldiv.quotient_msk\[5\] _2173_ _2156_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__mux2_1
X_4688_ _2110_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__inv_2
X_3708_ u_bits.i_op2\[9\] _1250_ _1272_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__a21oi_1
X_3639_ _0454_ _1368_ _1370_ _1371_ _1357_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__o221a_1
X_5309_ u_muldiv.divisor\[21\] _2616_ _2617_ u_muldiv.divisor\[22\] vssd1 vssd1 vccd1
+ vccd1 _0412_ sky130_fd_sc_hd__a22o_1
X_3990_ _1641_ _1648_ _1649_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__a21o_1
X_2941_ _0752_ _0753_ _0648_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__mux2_1
X_5660_ clknet_leaf_27_i_clk _0303_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[6\] sky130_fd_sc_hd__dfxtp_1
X_4611_ u_muldiv.dividend\[21\] u_muldiv.divisor\[21\] vssd1 vssd1 vccd1 vccd1 _2034_
+ sky130_fd_sc_hd__and2b_1
X_2872_ _0642_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__buf_2
X_5591_ clknet_leaf_37_i_clk _0238_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[8\] sky130_fd_sc_hd__dfxtp_1
X_4542_ u_muldiv.mul\[30\] o_add[0] _1583_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__mux2_1
X_4473_ u_bits.i_op2\[30\] _1966_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__xnor2_1
X_3424_ _1171_ _1194_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__xnor2_1
X_3355_ _0561_ _1138_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__xor2_4
X_3286_ _0788_ _1080_ _0911_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__o21a_1
X_5025_ u_muldiv.dividend\[8\] _2377_ _2378_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__mux2_1
X_4809_ u_muldiv.o_div\[15\] _2210_ u_muldiv.o_div\[16\] vssd1 vssd1 vccd1 vccd1 _2217_
+ sky130_fd_sc_hd__o21ai_1
X_5789_ clknet_leaf_38_i_clk _0431_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[37\] sky130_fd_sc_hd__dfxtp_1
X_3140_ _0944_ _0870_ _0774_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__mux2_1
X_3071_ u_bits.i_op1\[7\] u_bits.i_op1\[6\] u_bits.i_op1\[5\] u_bits.i_op1\[4\] _0657_
+ _0648_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__mux4_2
X_5712_ clknet_leaf_32_i_clk _0355_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_3973_ _1634_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__buf_2
X_2924_ _0467_ _0468_ _0737_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__a21bo_1
X_2855_ _0524_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__buf_4
X_5643_ clknet_leaf_40_i_clk _0290_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_5574_ clknet_leaf_9_i_clk _0221_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_4525_ _1994_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__clkbuf_1
X_2786_ _0568_ _0576_ _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__a21o_1
X_4456_ _1832_ _1953_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__nor2_1
X_3407_ o_add[0] o_add[1] vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__nor2_1
X_4387_ u_muldiv.divisor\[43\] _1867_ _1887_ u_muldiv.divisor\[44\] _1898_ vssd1 vssd1
+ vccd1 vccd1 _0209_ sky130_fd_sc_hd__a221o_1
X_3338_ _0532_ _0544_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__nand2_1
X_3269_ _1050_ _1065_ _0447_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__a21o_1
X_5008_ u_bits.i_op1\[4\] u_bits.i_op1\[5\] u_bits.i_op1\[6\] _2328_ vssd1 vssd1 vccd1
+ vccd1 _2363_ sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_31_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_46_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2640_ u_muldiv.i_op2_signed alu_ctrl\[2\] vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__nor2_4
X_5290_ _1209_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__buf_2
X_4310_ u_muldiv.divisor\[31\] vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__inv_2
X_4241_ _1794_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
X_4172_ o_wdata[4] i_reg_data2[4] _1756_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__mux2_1
X_3123_ _0908_ _0913_ _0929_ _0747_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__o31a_1
X_3054_ _0861_ _0862_ _0696_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__mux2_1
X_3956_ _1630_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__clkbuf_1
X_2907_ _0619_ _0625_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__nor2_2
X_3887_ _1214_ _1591_ _1592_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__and3_1
X_5626_ clknet_leaf_43_i_clk _0273_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_2838_ u_bits.i_op1\[16\] vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__buf_4
X_5557_ clknet_leaf_7_i_clk _0204_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_2769_ _0582_ _0583_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__xor2_4
X_4508_ _1985_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
X_5488_ clknet_leaf_51_i_clk _0136_ vssd1 vssd1 vccd1 vccd1 o_wdata[6] sky130_fd_sc_hd__dfxtp_4
X_4439_ u_bits.i_op2\[23\] _1938_ vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__or2_1
X_4790_ u_muldiv.quotient_msk\[12\] u_muldiv.o_div\[12\] _1841_ vssd1 vssd1 vccd1
+ vccd1 _2202_ sky130_fd_sc_hd__o21a_1
X_3810_ _0618_ _0639_ _1530_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__and3_1
X_3741_ u_muldiv.mul\[11\] _1330_ _1400_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__o21ai_1
X_3672_ _1106_ csr_data\[6\] _1388_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__o21ai_1
X_5411_ clknet_leaf_49_i_clk _0059_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[2\] sky130_fd_sc_hd__dfxtp_2
X_5342_ _1145_ _2628_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__nor2_1
X_5273_ u_muldiv.dividend\[30\] _2157_ _2604_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__a21o_1
X_4224_ u_wr_mux.i_reg_data2\[29\] i_reg_data2[29] _1778_ vssd1 vssd1 vccd1 vccd1
+ _1786_ sky130_fd_sc_hd__mux2_1
X_4155_ _0454_ i_alu_ctrl[1] _1745_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__mux2_1
X_3106_ _0644_ _0912_ _0712_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__o21a_1
X_4086_ _1715_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__clkbuf_1
X_3037_ _0739_ csr_data\[22\] _0847_ _0732_ vssd1 vssd1 vccd1 vccd1 o_result[22] sky130_fd_sc_hd__o211a_2
X_4988_ _2344_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__clkbuf_1
X_3939_ _0691_ i_op1[22] _1621_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__mux2_1
X_5609_ clknet_leaf_33_i_clk _0256_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[26\] sky130_fd_sc_hd__dfxtp_1
X_4911_ _1946_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__buf_2
X_4842_ _2153_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__buf_4
X_4773_ u_muldiv.o_div\[8\] _2188_ _2154_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__mux2_1
X_3724_ _0714_ _1449_ _1450_ _0624_ _1151_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__o32a_1
X_3655_ _0454_ _1382_ _1385_ _1386_ _1357_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__o221a_1
X_3586_ _1265_ _1318_ _1320_ _0906_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__o211ai_1
X_5325_ u_muldiv.divisor\[0\] u_muldiv.dividend\[0\] vssd1 vssd1 vccd1 vccd1 _2622_
+ sky130_fd_sc_hd__or2b_1
X_5256_ _0697_ _2588_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__xnor2_1
X_4207_ u_wr_mux.i_reg_data2\[21\] i_reg_data2[21] _1767_ vssd1 vssd1 vccd1 vccd1
+ _1777_ sky130_fd_sc_hd__mux2_1
X_5187_ u_muldiv.dividend\[22\] _2506_ u_muldiv.dividend\[23\] vssd1 vssd1 vccd1 vccd1
+ _2526_ sky130_fd_sc_hd__o21ai_1
X_4138_ o_pc_target[12] i_pc_target[12] _1734_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__mux2_1
X_4069_ u_bits.i_op2\[28\] _1687_ _1596_ i_op2[28] vssd1 vssd1 vccd1 vccd1 _1705_
+ sky130_fd_sc_hd__a22o_1
X_3440_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__clkbuf_4
X_3371_ _1152_ _0607_ _0578_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__a21o_1
X_5110_ _2456_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__clkbuf_1
X_5041_ u_muldiv.dividend\[10\] _2380_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__xor2_1
X_4825_ u_muldiv.quotient_msk\[19\] _2226_ _2229_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__mux2_1
X_4756_ _2165_ u_muldiv.o_div\[5\] _2173_ _1913_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__a31o_1
X_4687_ u_muldiv.divisor\[24\] u_muldiv.dividend\[24\] vssd1 vssd1 vccd1 vccd1 _2110_
+ sky130_fd_sc_hd__xor2_1
X_3707_ _0908_ _1434_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__nor2_1
X_3638_ u_muldiv.mul\[4\] _1330_ _1331_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__o21ai_1
X_3569_ _1124_ u_pc_sel.i_pc_next\[1\] _1304_ vssd1 vssd1 vccd1 vccd1 o_result[1]
+ sky130_fd_sc_hd__o21a_2
X_5308_ u_muldiv.divisor\[20\] _2616_ _2617_ u_muldiv.divisor\[21\] vssd1 vssd1 vccd1
+ vccd1 _0411_ sky130_fd_sc_hd__a22o_1
X_5239_ u_muldiv.dividend\[27\] _2164_ _2573_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__o21a_1
X_2940_ u_bits.i_op1\[23\] u_bits.i_op1\[24\] _0649_ vssd1 vssd1 vccd1 vccd1 _0753_
+ sky130_fd_sc_hd__mux2_1
X_2871_ _0634_ _0641_ _0685_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__and3_1
X_4610_ u_muldiv.divisor\[20\] u_muldiv.dividend\[20\] vssd1 vssd1 vccd1 vccd1 _2033_
+ sky130_fd_sc_hd__or2b_1
X_5590_ clknet_leaf_24_i_clk _0237_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[7\] sky130_fd_sc_hd__dfxtp_1
X_4541_ _2002_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__clkbuf_1
X_4472_ u_bits.i_op2\[29\] _1962_ _1845_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__o21a_1
X_3423_ _1070_ _1094_ _1101_ _1193_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__a31oi_4
X_3354_ _1141_ vssd1 vssd1 vccd1 vccd1 o_add[7] sky130_fd_sc_hd__inv_2
X_3285_ _0758_ _0823_ _0704_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__o21a_1
X_5024_ _2153_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__buf_4
X_4808_ _2181_ _2214_ _2216_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__a21oi_1
X_5788_ clknet_leaf_38_i_clk _0430_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[36\] sky130_fd_sc_hd__dfxtp_1
X_4739_ _2153_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__clkbuf_4
X_3070_ _0673_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__buf_4
X_5711_ clknet_leaf_33_i_clk _0354_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_3972_ i_inst_branch _1632_ _1636_ u_pc_sel.i_inst_branch vssd1 vssd1 vccd1 vccd1
+ _0056_ sky130_fd_sc_hd__a22o_1
X_2923_ _0470_ _0615_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__nand2_1
X_2854_ _0668_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__clkbuf_4
X_5642_ clknet_leaf_41_i_clk _0289_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_5573_ clknet_leaf_9_i_clk _0220_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_2785_ _0579_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__or2_1
X_4524_ u_muldiv.mul\[21\] u_muldiv.mul\[22\] _1989_ vssd1 vssd1 vccd1 vccd1 _1994_
+ sky130_fd_sc_hd__mux2_1
X_4455_ u_bits.i_op2\[26\] _1952_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__xnor2_1
X_3406_ _0538_ _0542_ vssd1 vssd1 vccd1 vccd1 o_add[1] sky130_fd_sc_hd__xor2_4
X_4386_ _1896_ _1897_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__nor2_1
X_3337_ _1128_ vssd1 vssd1 vccd1 vccd1 o_add[3] sky130_fd_sc_hd__inv_2
X_3268_ _0750_ o_add[29] _1063_ _1064_ _0804_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__a221o_1
X_5007_ _2293_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__buf_2
X_3199_ _0644_ _0999_ _0712_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__o21a_1
X_4240_ csr_data\[3\] i_csr_data[3] _1789_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__mux2_1
X_4171_ _1758_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__clkbuf_1
X_3122_ _0914_ _0921_ _0924_ _0925_ _0928_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__a221o_1
X_3053_ _0756_ _0761_ _0663_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__mux2_1
X_3955_ _0699_ i_op1[30] _1621_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__mux2_1
X_2906_ _0633_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__buf_2
X_5625_ clknet_leaf_43_i_clk _0272_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_3886_ u_muldiv.i_op2_signed _0626_ _1194_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__o21ai_1
X_2837_ _0630_ _0645_ _0646_ _0647_ _0648_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__mux4_1
X_5556_ clknet_leaf_7_i_clk _0203_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_2768_ u_bits.i_op1\[11\] u_muldiv.add_prev\[11\] _0450_ vssd1 vssd1 vccd1 vccd1
+ _0583_ sky130_fd_sc_hd__mux2_2
X_4507_ u_muldiv.mul\[13\] u_muldiv.mul\[14\] _1978_ vssd1 vssd1 vccd1 vccd1 _1985_
+ sky130_fd_sc_hd__mux2_1
X_2699_ u_bits.i_op1\[13\] u_muldiv.add_prev\[13\] _0449_ vssd1 vssd1 vccd1 vccd1
+ _0514_ sky130_fd_sc_hd__mux2_1
X_5487_ clknet_leaf_51_i_clk _0135_ vssd1 vssd1 vccd1 vccd1 o_wdata[5] sky130_fd_sc_hd__dfxtp_4
X_4438_ u_bits.i_op2\[23\] _1938_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__nand2_1
X_4369_ _1868_ _1883_ u_bits.i_op2\[9\] vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__a21oi_1
X_3740_ u_muldiv.mul\[43\] _1325_ _1465_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__a21oi_1
X_3671_ _0454_ _1397_ _1399_ _1401_ _1357_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__o221a_1
X_5410_ clknet_leaf_49_i_clk _0058_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[1\] sky130_fd_sc_hd__dfxtp_1
X_5341_ _1147_ _2628_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__nor2_1
X_5272_ _1209_ _2600_ _2603_ _2161_ vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__o211a_1
X_4223_ _1785_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__clkbuf_1
X_4154_ _1749_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__clkbuf_1
X_3105_ _0909_ _0910_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__o21a_1
X_4085_ u_pc_sel.i_pc_next\[3\] i_pc_next[3] _1712_ vssd1 vssd1 vccd1 vccd1 _1715_
+ sky130_fd_sc_hd__mux2_1
X_3036_ _0817_ _0846_ _0447_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_30_i_clk clknet_2_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4987_ u_muldiv.dividend\[5\] _2343_ _2244_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__mux2_1
X_3938_ _1595_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__clkbuf_4
X_3869_ _1583_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_45_i_clk clknet_2_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5608_ clknet_leaf_33_i_clk _0255_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[25\] sky130_fd_sc_hd__dfxtp_1
X_5539_ clknet_leaf_15_i_clk _0187_ vssd1 vssd1 vccd1 vccd1 csr_data\[23\] sky130_fd_sc_hd__dfxtp_1
X_4910_ u_muldiv.quotient_msk\[19\] _2282_ _2281_ u_muldiv.quotient_msk\[20\] vssd1
+ vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__a22o_1
X_4841_ _2208_ _2240_ _2241_ _2242_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__a31o_1
X_4772_ _1835_ _2185_ _2186_ _2187_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__a31o_1
X_3723_ _1445_ _1305_ _1272_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__a21oi_1
X_3654_ u_muldiv.mul\[5\] _1330_ _1331_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__o21ai_1
X_3585_ _0923_ _1255_ _1293_ _1319_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__a2bb2o_1
X_5324_ _1913_ _2621_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__nor2_1
X_5255_ _0996_ _1029_ _2568_ _2292_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__o31a_1
X_4206_ _1776_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__clkbuf_1
X_5186_ u_muldiv.dividend\[23\] u_muldiv.dividend\[22\] _2506_ vssd1 vssd1 vccd1 vccd1
+ _2525_ sky130_fd_sc_hd__or3_1
X_4137_ _1740_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__clkbuf_1
X_4068_ u_bits.i_op2\[29\] u_bits.i_op2\[27\] _1198_ vssd1 vssd1 vccd1 vccd1 _1704_
+ sky130_fd_sc_hd__mux2_1
X_3019_ _0691_ u_bits.i_op2\[22\] _0637_ _0829_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__o22a_1
X_3370_ _0568_ _0576_ _0599_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__a21o_1
X_5040_ _2392_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__clkbuf_1
X_4824_ _1206_ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__buf_4
X_4755_ u_muldiv.o_div\[4\] _2171_ _2174_ _2164_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__a22o_1
X_3706_ _1110_ _0949_ _1431_ _1249_ _1433_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__a221o_1
X_4686_ _2107_ _2108_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__nor2_1
X_3637_ u_muldiv.mul\[36\] _1325_ _1369_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__a21oi_1
X_3568_ _0446_ csr_data\[1\] _1300_ _1303_ _0730_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__a221o_1
X_5307_ u_muldiv.divisor\[19\] _2616_ _2617_ u_muldiv.divisor\[20\] vssd1 vssd1 vccd1
+ vccd1 _0410_ sky130_fd_sc_hd__a22o_1
X_3499_ o_wdata[7] _1233_ _0799_ u_wr_mux.i_reg_data2\[15\] vssd1 vssd1 vccd1 vccd1
+ _1241_ sky130_fd_sc_hd__a22o_1
X_5238_ _1209_ _2564_ _2565_ _2157_ _2572_ vssd1 vssd1 vccd1 vccd1 _2573_ sky130_fd_sc_hd__a311o_1
X_5169_ _2508_ _2509_ vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__xnor2_1
X_2870_ _0644_ _0671_ _0684_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__o21ai_1
X_4540_ u_muldiv.mul\[29\] u_muldiv.mul\[30\] _1583_ vssd1 vssd1 vccd1 vccd1 _2002_
+ sky130_fd_sc_hd__mux2_1
X_4471_ u_muldiv.divisor\[60\] _1836_ _1946_ u_muldiv.divisor\[61\] _1965_ vssd1 vssd1
+ vccd1 vccd1 _0226_ sky130_fd_sc_hd__a221o_1
X_3422_ _1102_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__inv_2
X_3353_ _0556_ _1140_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__xnor2_4
X_3284_ u_muldiv.mul\[30\] _0740_ _0720_ u_muldiv.mul\[62\] _1078_ vssd1 vssd1 vccd1
+ vccd1 _1079_ sky130_fd_sc_hd__a221o_1
X_5023_ _1878_ _2369_ _2376_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__o21a_1
X_4807_ _2167_ _2215_ u_muldiv.o_div\[15\] vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__a21oi_1
X_5787_ clknet_leaf_38_i_clk _0429_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[35\] sky130_fd_sc_hd__dfxtp_1
X_2999_ _0808_ _0809_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__or2_1
X_4738_ _1209_ _2158_ _2159_ _1842_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__a31o_1
X_4669_ _2090_ _2091_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__and2b_1
X_3971_ i_inst_jal_jalr _1632_ _1636_ u_pc_sel.i_inst_jal_jalr vssd1 vssd1 vccd1 vccd1
+ _0055_ sky130_fd_sc_hd__a22o_1
X_5710_ clknet_leaf_33_i_clk _0353_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_2922_ _0734_ _0735_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__xnor2_4
X_2853_ u_bits.i_op2\[2\] vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__clkbuf_4
X_5641_ clknet_leaf_40_i_clk _0288_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_2784_ _0590_ _0594_ _0598_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__or3_1
X_5572_ clknet_leaf_2_i_clk _0219_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_4523_ _1993_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__clkbuf_1
X_4454_ _1942_ _1951_ _1845_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__o21a_1
X_3405_ _0541_ _0540_ vssd1 vssd1 vccd1 vccd1 o_add[0] sky130_fd_sc_hd__xor2_4
X_4385_ u_bits.i_op2\[12\] _1852_ _1895_ _1856_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__a31o_1
X_3336_ _1126_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__xnor2_4
X_5006_ u_muldiv.dividend\[7\] _2345_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__or2_1
X_3267_ _0629_ _1059_ _0955_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__a21oi_1
X_3198_ _0909_ _0998_ _0911_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__o21a_1
X_4170_ o_wdata[3] i_reg_data2[3] _1756_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__mux2_1
X_3121_ _0904_ _0905_ _0926_ _0927_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__o22a_1
X_3052_ _0753_ _0755_ _0663_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__mux2_1
X_3954_ _1629_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__clkbuf_1
X_2905_ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__buf_2
X_3885_ u_muldiv.i_op2_signed _0626_ _1194_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__or3_1
X_5624_ clknet_leaf_44_i_clk _0271_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2836_ _0650_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__buf_4
X_5555_ clknet_leaf_8_i_clk _0202_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_2767_ _0456_ _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__xnor2_4
X_4506_ _1984_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
X_2698_ _0456_ _0512_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__xnor2_1
X_5486_ clknet_leaf_51_i_clk _0134_ vssd1 vssd1 vccd1 vccd1 o_wdata[4] sky130_fd_sc_hd__dfxtp_4
X_4437_ u_bits.i_op2\[22\] _1934_ _1846_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__o21ai_1
X_4368_ _1406_ u_bits.i_op2\[8\] _1873_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__or3_1
X_4299_ _1824_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
X_3319_ _0783_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__buf_4
X_3670_ u_muldiv.mul\[6\] _1330_ _1400_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__o21ai_1
X_5340_ _1584_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__buf_2
X_5271_ _2601_ _2602_ _1835_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__o21ai_1
X_4222_ u_wr_mux.i_reg_data2\[28\] i_reg_data2[28] _1778_ vssd1 vssd1 vccd1 vccd1
+ _1785_ sky130_fd_sc_hd__mux2_1
X_4153_ _1639_ i_alu_ctrl[0] _1745_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__mux2_1
X_3104_ _0524_ _0703_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__nand2_4
X_4084_ _1714_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__clkbuf_1
X_3035_ _0750_ o_add[22] _0844_ _0845_ _0804_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__a221o_1
X_4986_ _2208_ _2335_ _2336_ _2342_ vssd1 vssd1 vccd1 vccd1 _2343_ sky130_fd_sc_hd__a31o_1
X_3937_ _1620_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__clkbuf_1
X_3868_ _1582_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__buf_2
X_3799_ u_muldiv.dividend\[15\] _0742_ _0743_ u_muldiv.o_div\[15\] _0622_ vssd1 vssd1
+ vccd1 vccd1 _1521_ sky130_fd_sc_hd__a221o_1
X_5607_ clknet_leaf_33_i_clk _0254_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[24\] sky130_fd_sc_hd__dfxtp_1
X_2819_ _0620_ _0633_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__nand2_2
X_5538_ clknet_leaf_15_i_clk _0186_ vssd1 vssd1 vccd1 vccd1 csr_data\[22\] sky130_fd_sc_hd__dfxtp_1
X_5469_ clknet_leaf_13_i_clk _0117_ vssd1 vssd1 vccd1 vccd1 o_pc_target[11] sky130_fd_sc_hd__dfxtp_2
X_4840_ u_muldiv.quotient_msk\[22\] u_muldiv.o_div\[22\] _1840_ vssd1 vssd1 vccd1
+ vccd1 _2242_ sky130_fd_sc_hd__o21a_1
X_4771_ u_muldiv.quotient_msk\[8\] u_muldiv.o_div\[8\] _1841_ vssd1 vssd1 vccd1 vccd1
+ _2187_ sky130_fd_sc_hd__o21a_1
X_3722_ _0908_ _1448_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__nor2_1
X_3653_ u_muldiv.mul\[37\] _1325_ _1384_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__a21oi_1
X_5323_ u_muldiv.quotient_msk\[0\] _2152_ u_muldiv.o_div\[0\] vssd1 vssd1 vccd1 vccd1
+ _2621_ sky130_fd_sc_hd__a21oi_1
X_3584_ _0923_ _1255_ _0867_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__a21o_1
X_5254_ _2030_ _2131_ _2585_ _1839_ vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__a31o_1
X_5185_ _2524_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__clkbuf_1
X_4205_ u_wr_mux.i_reg_data2\[20\] i_reg_data2[20] _1767_ vssd1 vssd1 vccd1 vccd1
+ _1776_ sky130_fd_sc_hd__mux2_1
X_4136_ o_pc_target[11] i_pc_target[11] _1734_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__mux2_1
X_4067_ _1689_ _1702_ _1703_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__a21o_1
X_3018_ _0618_ _0639_ _0828_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__and3_1
X_4969_ _2068_ _2058_ _2067_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_44_i_clk clknet_2_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4823_ _2170_ u_muldiv.o_div\[19\] _2226_ _2196_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__a31o_1
X_4754_ _2165_ _2172_ _2173_ _1842_ u_muldiv.quotient_msk\[4\] vssd1 vssd1 vccd1 vccd1
+ _2174_ sky130_fd_sc_hd__a32o_1
X_3705_ u_bits.i_op2\[9\] _1250_ _0926_ _1432_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__o22a_1
X_4685_ u_muldiv.dividend\[25\] u_muldiv.divisor\[25\] vssd1 vssd1 vccd1 vccd1 _2108_
+ sky130_fd_sc_hd__and2b_1
X_3636_ u_muldiv.dividend\[4\] _1326_ _1327_ u_muldiv.o_div\[4\] _0717_ vssd1 vssd1
+ vccd1 vccd1 _1369_ sky130_fd_sc_hd__a221o_1
X_3567_ _1301_ _1302_ _0728_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__o21a_1
X_5306_ _1842_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__buf_2
X_5237_ _2303_ _2567_ _2571_ vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__a21oi_1
X_3498_ _1192_ u_wr_mux.i_reg_data2\[30\] _1240_ vssd1 vssd1 vccd1 vccd1 o_wdata[30]
+ sky130_fd_sc_hd__a21o_2
X_5168_ _2499_ _2100_ _2033_ vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__o21ai_1
X_5099_ _2444_ _2445_ vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__nand2_1
X_4119_ o_pc_target[3] i_pc_target[3] _1723_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__mux2_1
X_4470_ _1963_ _1964_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__nor2_1
X_3421_ _0619_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__clkbuf_8
X_3352_ _0561_ _1139_ _0570_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__o21a_1
X_3283_ u_muldiv.dividend\[30\] _0721_ _0723_ u_muldiv.o_div\[30\] _0744_ vssd1 vssd1
+ vccd1 vccd1 _1078_ sky130_fd_sc_hd__a221o_1
X_5022_ _2371_ _2372_ _2374_ _2375_ _1207_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__a221o_1
X_4806_ u_muldiv.quotient_msk\[15\] _2210_ _2156_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__mux2_1
X_5786_ clknet_leaf_38_i_clk _0428_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[34\] sky130_fd_sc_hd__dfxtp_1
X_2998_ _0808_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__nand2_1
X_4737_ u_muldiv.o_div\[2\] _2026_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__nand2_1
X_4668_ u_muldiv.divisor\[17\] u_muldiv.dividend\[17\] vssd1 vssd1 vccd1 vccd1 _2091_
+ sky130_fd_sc_hd__or2b_1
X_3619_ _1274_ _1351_ _1352_ _0624_ _1128_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__o32a_1
X_4599_ _1204_ _2023_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__nor2_1
X_3970_ i_rd[4] _1632_ _1636_ o_rd[4] vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__a22o_1
X_2921_ u_bits.i_op1\[21\] u_muldiv.add_prev\[21\] _0451_ vssd1 vssd1 vccd1 vccd1
+ _0735_ sky130_fd_sc_hd__mux2_2
X_2852_ _0665_ _0666_ _0663_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__mux2_1
X_5640_ clknet_leaf_40_i_clk _0287_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_2783_ _0596_ _0597_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__xnor2_1
X_5571_ clknet_leaf_2_i_clk _0218_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_4522_ u_muldiv.mul\[20\] u_muldiv.mul\[21\] _1989_ vssd1 vssd1 vccd1 vccd1 _1993_
+ sky130_fd_sc_hd__mux2_1
X_4453_ _0905_ u_bits.i_op2\[25\] vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__or2_1
X_3404_ o_add[9] o_add[13] o_add[17] vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__or3_1
X_4384_ _1868_ _1895_ u_bits.i_op2\[12\] vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__a21oi_1
X_3335_ _0528_ _0545_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__and2b_1
X_3266_ _0628_ _1052_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__or3_1
X_5005_ u_muldiv.dividend\[7\] _2345_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__nand2_1
X_3197_ _0862_ _0859_ _0668_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__mux2_1
X_5769_ clknet_leaf_17_i_clk _0412_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_3120_ _0904_ _0905_ _0867_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__a21oi_1
X_3051_ _0704_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__and2_1
X_3953_ _0697_ i_op1[29] _1621_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__mux2_1
X_2904_ _0618_ _0718_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__nor2_1
X_3884_ _1590_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__clkbuf_1
X_5623_ clknet_leaf_44_i_clk _0270_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2835_ _0649_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__buf_4
X_5554_ clknet_leaf_8_i_clk _0201_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_2766_ _0449_ u_bits.i_op1\[11\] _0497_ _0580_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__a31o_1
X_4505_ u_muldiv.mul\[12\] u_muldiv.mul\[13\] _1978_ vssd1 vssd1 vccd1 vccd1 _1984_
+ sky130_fd_sc_hd__mux2_1
X_2697_ _0449_ u_bits.i_op1\[13\] _0497_ _0511_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__a31o_1
X_5485_ clknet_leaf_51_i_clk _0133_ vssd1 vssd1 vccd1 vccd1 o_wdata[3] sky130_fd_sc_hd__dfxtp_4
X_4436_ u_muldiv.divisor\[53\] _1878_ _1833_ _1936_ _1937_ vssd1 vssd1 vccd1 vccd1
+ _0219_ sky130_fd_sc_hd__o221a_1
X_4367_ u_muldiv.divisor\[39\] _1878_ _1829_ u_muldiv.divisor\[40\] _1882_ vssd1 vssd1
+ vccd1 vccd1 _0205_ sky130_fd_sc_hd__o221a_1
X_3318_ _0831_ _0699_ _0763_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__a21o_1
X_4298_ csr_data\[31\] i_csr_data[31] _1595_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__mux2_1
X_3249_ _1045_ _1046_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__or2_2
X_5270_ u_muldiv.dividend\[30\] _2583_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__and2_1
X_4221_ _1784_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__clkbuf_1
X_4152_ _1748_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__clkbuf_1
X_3103_ _0690_ _0701_ _0668_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__mux2_1
X_4083_ u_pc_sel.i_pc_next\[2\] i_pc_next[2] _1712_ vssd1 vssd1 vccd1 vccd1 _1714_
+ sky130_fd_sc_hd__mux2_1
X_3034_ _0629_ _0828_ _0714_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__a21oi_1
X_4985_ _2229_ _2341_ vssd1 vssd1 vccd1 vccd1 _2342_ sky130_fd_sc_hd__nor2_1
X_3936_ _0768_ i_op1[21] _1610_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__mux2_1
X_3867_ _1198_ u_muldiv.i_on_wait vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__or2_1
X_5606_ clknet_leaf_33_i_clk _0253_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[23\] sky130_fd_sc_hd__dfxtp_1
X_2818_ _0632_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__buf_2
X_3798_ _0714_ _1518_ _1519_ _0623_ _1162_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__o32a_1
X_5537_ clknet_leaf_15_i_clk _0185_ vssd1 vssd1 vccd1 vccd1 csr_data\[21\] sky130_fd_sc_hd__dfxtp_1
X_2749_ _0456_ _0563_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__xnor2_4
X_5468_ clknet_leaf_13_i_clk _0116_ vssd1 vssd1 vccd1 vccd1 o_pc_target[10] sky130_fd_sc_hd__dfxtp_2
X_5399_ clknet_leaf_53_i_clk _0047_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[31\] sky130_fd_sc_hd__dfxtp_1
X_4419_ u_bits.i_op2\[19\] _1923_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__nand2_1
X_4770_ u_muldiv.o_div\[7\] u_muldiv.o_div\[8\] _2179_ vssd1 vssd1 vccd1 vccd1 _2186_
+ sky130_fd_sc_hd__or3_2
X_3721_ _1110_ _0975_ _1444_ _1248_ _1447_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__a221o_1
X_3652_ u_muldiv.dividend\[5\] _1326_ _1327_ u_muldiv.o_div\[5\] _1383_ vssd1 vssd1
+ vccd1 vccd1 _1384_ sky130_fd_sc_hd__a221o_1
X_3583_ _0669_ _0788_ _0840_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__or3b_1
X_5322_ u_muldiv.outsign _1913_ _2620_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__o21a_1
X_5253_ _2030_ _2131_ _2585_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__a21oi_1
X_5184_ u_muldiv.dividend\[22\] _2523_ _2485_ vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__mux2_1
X_4204_ _1775_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__clkbuf_1
X_4135_ _1739_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__clkbuf_1
X_4066_ u_bits.i_op2\[27\] _1687_ _1596_ i_op2[27] vssd1 vssd1 vccd1 vccd1 _1703_
+ sky130_fd_sc_hd__a22o_1
X_3017_ _0691_ u_bits.i_op2\[22\] vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__nand2_1
X_4968_ _2068_ _2058_ _2067_ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__nand3_1
X_4899_ _1946_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__buf_2
X_3919_ _1611_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__clkbuf_1
X_4822_ u_muldiv.o_div\[18\] _2171_ _2227_ _2164_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a22o_1
X_4753_ u_muldiv.o_div\[3\] u_muldiv.o_div\[4\] _2158_ vssd1 vssd1 vccd1 vccd1 _2173_
+ sky130_fd_sc_hd__or3_2
X_3704_ u_bits.i_op2\[9\] _1250_ _1267_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__a21oi_1
X_4684_ u_muldiv.divisor\[25\] u_muldiv.dividend\[25\] vssd1 vssd1 vccd1 vccd1 _2107_
+ sky130_fd_sc_hd__and2b_1
X_3635_ _1274_ _1366_ _1367_ _0624_ _1137_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__o32a_1
X_3566_ u_muldiv.dividend\[1\] _0721_ _0723_ u_muldiv.o_div\[1\] _0724_ vssd1 vssd1
+ vccd1 vccd1 _1302_ sky130_fd_sc_hd__a221o_1
X_5305_ u_muldiv.divisor\[18\] _2616_ _2615_ u_muldiv.divisor\[19\] vssd1 vssd1 vccd1
+ vccd1 _0409_ sky130_fd_sc_hd__a22o_1
X_3497_ o_wdata[6] _1233_ _0799_ u_wr_mux.i_reg_data2\[14\] vssd1 vssd1 vccd1 vccd1
+ _1240_ sky130_fd_sc_hd__a22o_1
X_5236_ _1207_ _2569_ _2570_ _1829_ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__o31a_1
X_5167_ _2034_ _2032_ vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__and2b_1
X_5098_ u_muldiv.dividend\[14\] _2423_ u_muldiv.dividend\[15\] vssd1 vssd1 vccd1 vccd1
+ _2445_ sky130_fd_sc_hd__o21ai_1
X_4118_ _1730_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__clkbuf_1
X_4049_ _1689_ _1690_ _1691_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__a21o_1
X_3420_ _0618_ _1170_ _1189_ _1190_ _0619_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__a221o_1
X_3351_ _1138_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__inv_2
X_3282_ _1072_ _1077_ vssd1 vssd1 vccd1 vccd1 o_add[30] sky130_fd_sc_hd__xor2_4
X_5021_ _1839_ vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__clkbuf_4
X_4805_ _2170_ u_muldiv.o_div\[15\] _2210_ _2196_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__a31o_1
X_5785_ clknet_leaf_35_i_clk _0427_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[33\] sky130_fd_sc_hd__dfxtp_1
X_2997_ u_bits.i_op1\[22\] u_muldiv.add_prev\[22\] _0451_ vssd1 vssd1 vccd1 vccd1
+ _0809_ sky130_fd_sc_hd__mux2_1
X_4736_ u_muldiv.o_div\[2\] _2026_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__or2_2
X_4667_ u_muldiv.dividend\[17\] u_muldiv.divisor\[17\] vssd1 vssd1 vccd1 vccd1 _2090_
+ sky130_fd_sc_hd__and2b_1
X_3618_ _0909_ _0794_ _1272_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__a21oi_1
X_4598_ op_cnt\[3\] op_cnt\[4\] _2020_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__and3_1
X_3549_ _1281_ _1282_ _1283_ _1284_ _0760_ _0879_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__mux4_1
X_5219_ u_muldiv.dividend\[25\] _2164_ _2555_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_43_i_clk clknet_2_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2920_ _0458_ _0733_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__xnor2_4
X_2851_ u_bits.i_op1\[6\] u_bits.i_op1\[5\] _0649_ vssd1 vssd1 vccd1 vccd1 _0666_
+ sky130_fd_sc_hd__mux2_1
X_2782_ u_bits.i_op1\[8\] u_muldiv.add_prev\[8\] _0450_ vssd1 vssd1 vccd1 vccd1 _0597_
+ sky130_fd_sc_hd__mux2_1
X_5570_ clknet_leaf_2_i_clk _0217_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_4521_ _1992_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__clkbuf_1
X_4452_ u_muldiv.divisor\[56\] _1836_ _1946_ u_muldiv.divisor\[57\] _1950_ vssd1 vssd1
+ vccd1 vccd1 _0222_ sky130_fd_sc_hd__a221o_1
X_3403_ _1176_ vssd1 vssd1 vccd1 vccd1 o_add[17] sky130_fd_sc_hd__inv_2
X_4383_ _1445_ u_bits.i_op2\[11\] _1888_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__or3_1
X_3334_ _0546_ _1125_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__nand2_2
X_3265_ _0914_ _1055_ _1058_ _0925_ _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__a221o_1
X_5004_ _2356_ _2357_ _2358_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__a21oi_1
X_3196_ _0996_ u_bits.i_op2\[27\] _0906_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__a21o_1
X_5768_ clknet_leaf_16_i_clk _0411_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_4719_ u_muldiv.divisor\[55\] u_muldiv.divisor\[54\] u_muldiv.divisor\[53\] u_muldiv.divisor\[52\]
+ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__or4_1
X_5699_ clknet_leaf_29_i_clk _0342_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3050_ u_bits.i_sra _0675_ _0702_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__o21a_1
X_3952_ _1628_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__clkbuf_1
X_2903_ _0639_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__clkbuf_4
X_3883_ o_add[31] _1579_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__and2_1
X_5622_ clknet_leaf_44_i_clk _0269_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_2834_ u_bits.i_op2\[0\] vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__buf_4
X_5553_ clknet_leaf_8_i_clk _0200_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_4504_ _1983_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__clkbuf_1
X_2765_ _0448_ u_bits.i_op2\[11\] vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__and2b_1
X_2696_ _0448_ u_bits.i_op2\[13\] vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__and2b_1
X_5484_ clknet_leaf_51_i_clk _0132_ vssd1 vssd1 vccd1 vccd1 o_wdata[2] sky130_fd_sc_hd__dfxtp_4
X_4435_ u_muldiv.divisor\[54\] _1829_ vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__or2_1
X_4366_ u_bits.i_op2\[8\] _1879_ _1881_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__a21o_1
X_3317_ _0925_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__buf_2
X_4297_ _1823_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
X_3248_ _1043_ _1044_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__nor2_1
X_3179_ _0628_ _0972_ _0981_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__or3_2
X_4220_ u_wr_mux.i_reg_data2\[27\] i_reg_data2[27] _1778_ vssd1 vssd1 vccd1 vccd1
+ _1784_ sky130_fd_sc_hd__mux2_1
X_4151_ _0618_ i_funct3[2] _1745_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__mux2_1
X_3102_ _0788_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__buf_4
X_4082_ _1713_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__clkbuf_1
X_3033_ _0628_ _0827_ _0830_ _0843_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__or4_1
X_4984_ _2337_ _2338_ _2340_ _1826_ vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__o22a_1
X_3935_ _1619_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__clkbuf_1
X_5605_ clknet_leaf_33_i_clk _0252_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[22\] sky130_fd_sc_hd__dfxtp_1
X_3866_ _1581_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__clkbuf_1
X_2817_ _0619_ o_funct3[2] vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__and2_1
X_3797_ u_bits.i_op2\[15\] _0654_ _0906_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__a21oi_1
X_5536_ clknet_leaf_15_i_clk _0184_ vssd1 vssd1 vccd1 vccd1 csr_data\[20\] sky130_fd_sc_hd__dfxtp_1
X_2748_ _0459_ u_bits.i_op2\[5\] u_bits.i_op1\[5\] _0463_ vssd1 vssd1 vccd1 vccd1
+ _0563_ sky130_fd_sc_hd__a22o_1
X_5467_ clknet_leaf_13_i_clk _0115_ vssd1 vssd1 vccd1 vccd1 o_pc_target[9] sky130_fd_sc_hd__dfxtp_2
X_2679_ _0488_ _0492_ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__a21o_1
X_4418_ u_bits.i_op2\[18\] _1919_ _1846_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__o21ai_1
X_5398_ clknet_leaf_4_i_clk _0046_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[30\] sky130_fd_sc_hd__dfxtp_2
X_4349_ _1835_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__buf_2
X_3720_ _1445_ _1305_ _0926_ _1446_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__o22a_1
X_3651_ _0622_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__buf_2
X_3582_ _1313_ _1316_ _0644_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__mux2_1
X_5321_ _1233_ _1115_ _2618_ _2619_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__a31o_1
X_5252_ _2133_ _2132_ vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__and2b_1
X_5183_ _2521_ _2522_ _2229_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__mux2_1
X_4203_ u_wr_mux.i_reg_data2\[19\] i_reg_data2[19] _1767_ vssd1 vssd1 vccd1 vccd1
+ _1775_ sky130_fd_sc_hd__mux2_1
X_4134_ o_pc_target[10] i_pc_target[10] _1734_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__mux2_1
X_4065_ u_bits.i_op2\[28\] u_bits.i_op2\[26\] _1681_ vssd1 vssd1 vccd1 vccd1 _1702_
+ sky130_fd_sc_hd__mux2_1
X_3016_ _0751_ _0826_ _0712_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__o21a_1
X_4967_ _2325_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__clkbuf_1
X_4898_ u_muldiv.quotient_msk\[9\] _2280_ _2279_ u_muldiv.quotient_msk\[10\] vssd1
+ vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__a22o_1
X_3918_ _0777_ i_op1[12] _1610_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__mux2_1
X_3849_ u_muldiv.mul\[19\] _0717_ _0720_ u_muldiv.mul\[51\] _1566_ vssd1 vssd1 vccd1
+ vccd1 _1567_ sky130_fd_sc_hd__a221o_1
X_5519_ clknet_leaf_13_i_clk _0167_ vssd1 vssd1 vccd1 vccd1 csr_data\[3\] sky130_fd_sc_hd__dfxtp_1
X_4821_ _2165_ _2225_ _2226_ _1842_ u_muldiv.quotient_msk\[18\] vssd1 vssd1 vccd1
+ vccd1 _2227_ sky130_fd_sc_hd__a32o_1
X_4752_ u_muldiv.o_div\[3\] _2158_ u_muldiv.o_div\[4\] vssd1 vssd1 vccd1 vccd1 _2172_
+ sky130_fd_sc_hd__o21ai_1
X_4683_ u_muldiv.divisor\[23\] u_muldiv.dividend\[23\] vssd1 vssd1 vccd1 vccd1 _2106_
+ sky130_fd_sc_hd__and2b_1
X_3703_ _1430_ _1289_ _0940_ _0824_ _0670_ _0643_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__mux4_1
X_3634_ _0688_ _1310_ _1272_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__a21oi_1
X_3565_ u_muldiv.mul\[1\] _0622_ _0719_ u_muldiv.mul\[33\] vssd1 vssd1 vccd1 vccd1
+ _1301_ sky130_fd_sc_hd__a22o_1
X_5304_ u_muldiv.divisor\[17\] _2616_ _2615_ u_muldiv.divisor\[18\] vssd1 vssd1 vccd1
+ vccd1 _0408_ sky130_fd_sc_hd__a22o_1
X_3496_ _1192_ u_wr_mux.i_reg_data2\[29\] _1239_ vssd1 vssd1 vccd1 vccd1 o_wdata[29]
+ sky130_fd_sc_hd__a21o_2
X_5235_ _2362_ _2568_ _0996_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__a21oi_1
X_5166_ u_muldiv.dividend\[20\] _2487_ u_muldiv.dividend\[21\] vssd1 vssd1 vccd1 vccd1
+ _2507_ sky130_fd_sc_hd__o21ai_1
X_5097_ u_muldiv.dividend\[15\] u_muldiv.dividend\[14\] _2423_ vssd1 vssd1 vccd1 vccd1
+ _2444_ sky130_fd_sc_hd__or3_2
X_4117_ o_pc_target[2] i_pc_target[2] _1723_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__mux2_1
X_4048_ u_bits.i_op2\[21\] _1687_ _1675_ i_op2[21] vssd1 vssd1 vccd1 vccd1 _1691_
+ sky130_fd_sc_hd__a22o_1
X_3350_ _1133_ _0566_ _0574_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__o21ai_4
X_5020_ _0785_ _2373_ vssd1 vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__xnor2_1
X_3281_ _1073_ _1075_ _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__and3_1
X_4804_ _2213_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__clkbuf_1
X_5784_ clknet_leaf_34_i_clk _0426_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[32\] sky130_fd_sc_hd__dfxtp_1
X_4735_ u_muldiv.outsign _2156_ _2152_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__a21oi_4
X_2996_ _0457_ _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__xnor2_1
X_4666_ _2087_ _2088_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__nand2_1
X_4597_ op_cnt\[3\] _2020_ _2022_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__o21a_1
X_3617_ _1249_ _1346_ _1350_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__a21oi_1
X_3548_ _1257_ _0786_ u_bits.i_op1\[7\] _0785_ _0778_ _0783_ vssd1 vssd1 vccd1 vccd1
+ _1284_ sky130_fd_sc_hd__mux4_1
X_3479_ _1230_ vssd1 vssd1 vccd1 vccd1 o_wdata[21] sky130_fd_sc_hd__buf_2
X_5218_ _1829_ _2547_ _2554_ _2154_ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__o211a_1
X_5149_ u_bits.i_op1\[17\] u_bits.i_op1\[18\] _2469_ vssd1 vssd1 vccd1 vccd1 _2492_
+ sky130_fd_sc_hd__or3_2
X_2850_ u_bits.i_op1\[8\] u_bits.i_op1\[7\] _0649_ vssd1 vssd1 vccd1 vccd1 _0665_
+ sky130_fd_sc_hd__mux2_1
X_2781_ _0457_ _0595_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__xnor2_2
X_4520_ u_muldiv.mul\[20\] u_muldiv.mul\[19\] _1214_ vssd1 vssd1 vccd1 vccd1 _1992_
+ sky130_fd_sc_hd__mux2_1
X_4451_ _1948_ _1949_ _1833_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__a21oi_1
X_3402_ _0610_ _1175_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__xor2_2
X_4382_ u_muldiv.divisor\[42\] _1867_ _1887_ u_muldiv.divisor\[43\] _1894_ vssd1 vssd1
+ vccd1 vccd1 _0208_ sky130_fd_sc_hd__a221o_1
X_3333_ _0532_ _0544_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__or2_1
X_3264_ _0697_ u_bits.i_op2\[29\] _0636_ _1060_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__o22a_1
X_5003_ _2356_ _2357_ _1841_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__o21ai_1
X_3195_ u_bits.i_op1\[27\] vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__clkbuf_4
X_5767_ clknet_leaf_16_i_clk _0410_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_2979_ _0791_ u_bits.i_op1\[0\] _0650_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__mux2_1
X_5698_ clknet_leaf_29_i_clk _0341_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4718_ u_muldiv.divisor\[35\] u_muldiv.divisor\[34\] u_muldiv.divisor\[33\] u_muldiv.divisor\[32\]
+ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__or4_1
X_4649_ u_muldiv.dividend\[6\] u_muldiv.divisor\[6\] vssd1 vssd1 vccd1 vccd1 _2072_
+ sky130_fd_sc_hd__and2b_1
X_3951_ _1029_ i_op1[28] _1621_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__mux2_1
X_2902_ _0622_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__clkbuf_4
X_3882_ _1589_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__clkbuf_1
X_5621_ clknet_leaf_46_i_clk _0268_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2833_ _0533_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__clkbuf_4
X_5552_ clknet_leaf_8_i_clk _0199_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_2764_ _0510_ _0577_ _0578_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__or3_1
X_4503_ u_muldiv.mul\[11\] u_muldiv.mul\[12\] _1978_ vssd1 vssd1 vccd1 vccd1 _1983_
+ sky130_fd_sc_hd__mux2_1
X_2695_ _0508_ _0502_ _0509_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__or3_1
X_5483_ clknet_leaf_51_i_clk _0131_ vssd1 vssd1 vccd1 vccd1 o_wdata[1] sky130_fd_sc_hd__dfxtp_4
X_4434_ u_bits.i_op2\[22\] _1935_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__xnor2_1
X_4365_ u_bits.i_op2\[8\] _1879_ _1880_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__o21ai_1
X_3316_ _0877_ _0882_ _0670_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__mux2_1
X_4296_ csr_data\[30\] i_csr_data[30] _1595_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__mux2_1
X_3247_ _1043_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_42_i_clk clknet_2_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3178_ _0914_ _0975_ _0977_ _0925_ _0980_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__a221o_1
X_4150_ _1747_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__clkbuf_1
X_3101_ _0858_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__buf_2
X_4081_ u_pc_sel.i_pc_next\[1\] i_pc_next[1] _1712_ vssd1 vssd1 vccd1 vccd1 _1713_
+ sky130_fd_sc_hd__mux2_1
X_3032_ _0672_ _0837_ _0842_ _0800_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__o211a_1
X_4983_ _1257_ _2339_ vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__xnor2_1
X_3934_ _0630_ i_op1[20] _1610_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__mux2_1
X_3865_ o_add[22] _1579_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__and2_1
X_5604_ clknet_leaf_33_i_clk _0251_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[21\] sky130_fd_sc_hd__dfxtp_1
X_2816_ _0630_ u_bits.i_op2\[20\] vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__nand2_1
X_3796_ _1514_ _1517_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__nor2_1
X_5535_ clknet_leaf_16_i_clk _0183_ vssd1 vssd1 vccd1 vccd1 csr_data\[19\] sky130_fd_sc_hd__dfxtp_1
X_2747_ _0556_ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__or2_1
X_5466_ clknet_leaf_13_i_clk _0114_ vssd1 vssd1 vccd1 vccd1 o_pc_target[8] sky130_fd_sc_hd__dfxtp_2
X_2678_ _0486_ _0487_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__nor2_1
X_4417_ u_muldiv.divisor\[49\] _1878_ _1833_ _1921_ _1922_ vssd1 vssd1 vccd1 vccd1
+ _0215_ sky130_fd_sc_hd__o221a_1
X_5397_ clknet_leaf_4_i_clk _0045_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[29\] sky130_fd_sc_hd__dfxtp_1
X_4348_ u_muldiv.divisor\[36\] _1838_ _1843_ u_muldiv.divisor\[37\] _1866_ vssd1 vssd1
+ vccd1 vccd1 _0202_ sky130_fd_sc_hd__a221o_1
X_4279_ _1814_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__clkbuf_1
X_3650_ _1274_ _1380_ _1381_ _0624_ _1135_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__o32a_1
X_3581_ _0970_ _1315_ _0879_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__mux2_1
X_5320_ _0619_ _2362_ _1831_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__a21o_1
X_5251_ u_muldiv.dividend\[28\] _2564_ u_muldiv.dividend\[29\] vssd1 vssd1 vccd1 vccd1
+ _2584_ sky130_fd_sc_hd__o21ai_1
X_4202_ _1774_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__clkbuf_1
X_5182_ u_muldiv.dividend\[22\] _2506_ vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__xor2_1
X_4133_ _1738_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__clkbuf_1
X_4064_ _1689_ _1700_ _1701_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__a21o_1
X_3015_ _0818_ _0822_ _0823_ _0824_ _0825_ _0707_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__mux4_2
X_4966_ u_muldiv.dividend\[3\] _2324_ _2244_ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__mux2_1
X_4897_ u_muldiv.quotient_msk\[8\] _2280_ _2279_ u_muldiv.quotient_msk\[9\] vssd1
+ vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__a22o_1
X_3917_ _1595_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__clkbuf_4
X_3848_ u_muldiv.dividend\[19\] _0721_ _0723_ u_muldiv.o_div\[19\] _0724_ vssd1 vssd1
+ vccd1 vccd1 _1566_ sky130_fd_sc_hd__a221o_1
X_3779_ u_bits.i_op2\[14\] _0655_ _0926_ _1501_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__o22a_1
X_5518_ clknet_leaf_13_i_clk _0166_ vssd1 vssd1 vccd1 vccd1 csr_data\[2\] sky130_fd_sc_hd__dfxtp_1
X_5449_ clknet_leaf_2_i_clk _0097_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_4820_ u_muldiv.o_div\[17\] u_muldiv.o_div\[18\] _2218_ vssd1 vssd1 vccd1 vccd1 _2226_
+ sky130_fd_sc_hd__or3_2
X_4751_ u_muldiv.outsign _2170_ _1913_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__a21oi_4
X_4682_ _2035_ _2102_ _2104_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__a21oi_1
X_3702_ _1281_ _1282_ _0760_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__mux2_1
X_3633_ _1265_ _0681_ _1362_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__o211a_1
X_3564_ _1298_ _1299_ _0804_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__a21o_1
X_5303_ u_muldiv.divisor\[16\] _2616_ _2615_ u_muldiv.divisor\[17\] vssd1 vssd1 vccd1
+ vccd1 _0407_ sky130_fd_sc_hd__a22o_1
X_3495_ o_wdata[5] _1233_ _0799_ u_wr_mux.i_reg_data2\[13\] vssd1 vssd1 vccd1 vccd1
+ _1239_ sky130_fd_sc_hd__a22o_1
X_5234_ _0996_ _2295_ _2568_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__and3_1
X_5165_ u_muldiv.dividend\[21\] u_muldiv.dividend\[20\] _2487_ vssd1 vssd1 vccd1 vccd1
+ _2506_ sky130_fd_sc_hd__or3_1
X_4116_ _1729_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__clkbuf_1
X_5096_ _2443_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__clkbuf_1
X_4047_ u_bits.i_op2\[22\] u_bits.i_op2\[20\] _1681_ vssd1 vssd1 vccd1 vccd1 _1690_
+ sky130_fd_sc_hd__mux2_1
X_4949_ _1255_ _2293_ _2308_ vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__and3_1
X_3280_ _1021_ _1046_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__or2_1
X_4803_ u_muldiv.o_div\[14\] _2212_ _2154_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__mux2_1
X_5783_ clknet_leaf_34_i_clk _0425_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[31\] sky130_fd_sc_hd__dfxtp_1
X_4734_ _1206_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__buf_4
X_2995_ _0460_ u_bits.i_op2\[22\] _0464_ u_bits.i_op1\[22\] vssd1 vssd1 vccd1 vccd1
+ _0807_ sky130_fd_sc_hd__a22o_1
X_4665_ u_muldiv.dividend\[16\] u_muldiv.divisor\[16\] vssd1 vssd1 vccd1 vccd1 _2088_
+ sky130_fd_sc_hd__or2b_1
X_4596_ _1204_ _2021_ vssd1 vssd1 vccd1 vccd1 _2022_ sky130_fd_sc_hd__nor2_1
X_3616_ _1265_ _1347_ _1349_ _0634_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__o211ai_1
X_3547_ _0791_ _1255_ _0794_ u_bits.i_op1\[4\] _0651_ _0783_ vssd1 vssd1 vccd1 vccd1
+ _1283_ sky130_fd_sc_hd__mux4_1
X_3478_ o_wdata[5] u_wr_mux.i_reg_data2\[21\] _1224_ vssd1 vssd1 vccd1 vccd1 _1230_
+ sky130_fd_sc_hd__mux2_1
X_5217_ _1831_ _2549_ _2550_ _2553_ _1877_ vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__o32a_1
X_5148_ _2094_ _2489_ _2490_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__a21o_1
X_5079_ u_bits.i_op1\[10\] u_bits.i_op1\[11\] u_bits.i_op1\[12\] _2394_ vssd1 vssd1
+ vccd1 vccd1 _2428_ sky130_fd_sc_hd__or4_4
X_2780_ _0460_ u_bits.i_op2\[8\] u_bits.i_op1\[8\] _0464_ vssd1 vssd1 vccd1 vccd1
+ _0595_ sky130_fd_sc_hd__a22o_1
X_4450_ u_bits.i_op2\[25\] _1947_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__or2_1
X_3401_ _0492_ _1164_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nand2_1
X_4381_ _1832_ _1893_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__nor2_1
X_3332_ _1106_ csr_data\[31\] _1123_ _1124_ vssd1 vssd1 vccd1 vccd1 o_result[31] sky130_fd_sc_hd__o211a_2
X_3263_ _0617_ _0638_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__and3_1
X_5002_ _2073_ _2055_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__nor2_1
X_3194_ u_muldiv.mul\[27\] _0740_ _0741_ u_muldiv.mul\[59\] _0994_ vssd1 vssd1 vccd1
+ vccd1 _0995_ sky130_fd_sc_hd__a221o_1
X_5766_ clknet_leaf_16_i_clk _0409_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_2978_ u_bits.i_op1\[1\] vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__clkbuf_4
X_5697_ clknet_leaf_29_i_clk _0340_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4717_ u_muldiv.divisor\[43\] u_muldiv.divisor\[42\] u_muldiv.divisor\[41\] _2139_
+ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__or4_1
X_4648_ _2057_ _2069_ _2070_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__o21ba_1
X_4579_ o_add[26] _2004_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__and2_1
X_3950_ _1627_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__clkbuf_1
X_2901_ _0616_ _0624_ _0715_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__o21ai_1
X_3881_ o_add[30] _1579_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__and2_1
X_5620_ clknet_leaf_46_i_clk _0267_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2832_ u_bits.i_op1\[17\] vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__buf_4
X_5551_ clknet_leaf_8_i_clk _0198_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_2763_ _0517_ _0518_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__xnor2_1
X_4502_ _1982_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__clkbuf_1
X_5482_ clknet_leaf_51_i_clk _0130_ vssd1 vssd1 vccd1 vccd1 o_wdata[0] sky130_fd_sc_hd__dfxtp_4
X_2694_ _0505_ _0506_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__xnor2_4
X_4433_ _1850_ _1934_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__nand2_1
X_4364_ u_muldiv.on_wait u_muldiv.i_on_end vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__nor2_4
X_4295_ _1822_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
X_3315_ u_muldiv.mul\[31\] _0740_ _0720_ u_muldiv.mul\[63\] _1107_ vssd1 vssd1 vccd1
+ vccd1 _1108_ sky130_fd_sc_hd__a221o_1
X_3246_ _0697_ u_muldiv.add_prev\[29\] _0452_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__mux2_1
X_3177_ _0689_ u_bits.i_op2\[26\] _0636_ _0979_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__o22a_1
X_5749_ clknet_leaf_24_i_clk _0392_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3100_ _0904_ _0905_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__a21o_1
X_4080_ _1711_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__clkbuf_4
X_3031_ _0674_ _0841_ _0642_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__a21bo_1
X_4982_ _1310_ _2328_ _2292_ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__o21a_1
X_3933_ _1618_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__clkbuf_1
X_3864_ _1580_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__clkbuf_1
X_5603_ clknet_leaf_33_i_clk _0250_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[20\] sky130_fd_sc_hd__dfxtp_1
X_2815_ u_bits.i_op1\[20\] vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__buf_4
X_3795_ _1110_ _1109_ _1516_ _0858_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__a211o_1
X_5534_ clknet_leaf_14_i_clk _0182_ vssd1 vssd1 vccd1 vccd1 csr_data\[18\] sky130_fd_sc_hd__dfxtp_1
X_2746_ _0559_ _0560_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__xnor2_4
X_5465_ clknet_leaf_13_i_clk _0113_ vssd1 vssd1 vccd1 vccd1 o_pc_target[7] sky130_fd_sc_hd__dfxtp_2
X_2677_ _0490_ _0491_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__nand2_1
X_4416_ u_muldiv.divisor\[50\] _1829_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__or2_1
X_5396_ clknet_leaf_4_i_clk _0044_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[28\] sky130_fd_sc_hd__dfxtp_2
X_4347_ _1864_ _1865_ _1833_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__a21oi_1
X_4278_ csr_data\[21\] i_csr_data[21] _1811_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__mux2_1
X_3229_ _0687_ _1027_ _0711_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__o21a_1
X_3580_ _1314_ _0818_ _0758_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_41_i_clk clknet_2_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5250_ u_muldiv.dividend\[29\] u_muldiv.dividend\[28\] _2564_ vssd1 vssd1 vccd1 vccd1
+ _2583_ sky130_fd_sc_hd__or3_1
X_4201_ u_wr_mux.i_reg_data2\[18\] i_reg_data2[18] _1767_ vssd1 vssd1 vccd1 vccd1
+ _1774_ sky130_fd_sc_hd__mux2_1
X_5181_ _2105_ _2518_ _2520_ _2375_ vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__a2bb2o_1
X_4132_ o_pc_target[9] i_pc_target[9] _1734_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__mux2_1
X_4063_ u_bits.i_op2\[26\] _1687_ _1596_ i_op2[26] vssd1 vssd1 vccd1 vccd1 _1701_
+ sky130_fd_sc_hd__a22o_1
X_3014_ _0696_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__buf_4
X_4965_ _2208_ _2315_ _2316_ _2323_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__a31o_1
X_3916_ _1609_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__clkbuf_1
X_4896_ u_muldiv.quotient_msk\[7\] _2280_ _2279_ u_muldiv.quotient_msk\[8\] vssd1
+ vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__a22o_1
X_3847_ _1106_ csr_data\[18\] _1565_ _1124_ vssd1 vssd1 vccd1 vccd1 o_result[18] sky130_fd_sc_hd__o211a_2
X_3778_ u_bits.i_op2\[14\] _0655_ _1267_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__a21oi_1
X_5517_ clknet_leaf_13_i_clk _0165_ vssd1 vssd1 vccd1 vccd1 csr_data\[1\] sky130_fd_sc_hd__dfxtp_1
X_2729_ _0538_ _0542_ _0543_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__a21oi_1
X_5448_ clknet_leaf_9_i_clk _0096_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_5379_ clknet_leaf_47_i_clk _0027_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[11\] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_2_0__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4750_ _2156_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__clkbuf_4
X_4681_ _2031_ _2103_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__or2_1
X_3701_ _1428_ _1429_ _1336_ u_pc_sel.i_pc_next\[8\] vssd1 vssd1 vccd1 vccd1 o_result[8]
+ sky130_fd_sc_hd__a2bb2o_2
X_3632_ _0858_ _1364_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__nor2_1
X_5302_ _1209_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__buf_2
X_3563_ _1112_ _0791_ _0906_ _0955_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__a211o_1
X_3494_ _1192_ u_wr_mux.i_reg_data2\[28\] _1238_ vssd1 vssd1 vccd1 vccd1 o_wdata[28]
+ sky130_fd_sc_hd__a21o_2
X_5233_ _0943_ _0689_ _2548_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__or3_1
X_5164_ _2505_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__clkbuf_1
X_4115_ o_pc_target[1] i_pc_target[1] _1723_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__mux2_1
X_5095_ u_muldiv.dividend\[14\] _2442_ _2378_ vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__mux2_1
X_4046_ _1635_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__buf_2
X_4948_ u_bits.i_op1\[0\] u_bits.i_op1\[1\] vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__or2_2
X_4879_ u_muldiv.quotient_msk\[30\] u_muldiv.o_div\[30\] vssd1 vssd1 vccd1 vccd1 _2273_
+ sky130_fd_sc_hd__or2_1
X_4802_ _2208_ _2209_ _2210_ _2211_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__a31o_1
X_5782_ clknet_leaf_24_i_clk _0424_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2994_ _0739_ csr_data\[21\] _0806_ _0732_ vssd1 vssd1 vccd1 vccd1 o_result[21] sky130_fd_sc_hd__o211a_2
X_4733_ _2155_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__clkbuf_1
X_4664_ u_muldiv.divisor\[16\] u_muldiv.dividend\[16\] vssd1 vssd1 vccd1 vccd1 _2087_
+ sky130_fd_sc_hd__or2b_1
X_4595_ op_cnt\[3\] _2020_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__and2_1
X_3615_ _0909_ _0794_ _1293_ _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__a2bb2o_1
X_3546_ u_bits.i_op1\[13\] _0655_ _0654_ _0653_ _0658_ _0779_ vssd1 vssd1 vccd1 vccd1
+ _1282_ sky130_fd_sc_hd__mux4_2
X_5216_ _2551_ _2552_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__nand2_1
X_3477_ _1229_ vssd1 vssd1 vccd1 vccd1 o_wdata[20] sky130_fd_sc_hd__buf_2
X_5147_ _2094_ _2489_ _1826_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__o21ai_1
X_5078_ _2044_ _2415_ _2425_ _2288_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__a31o_1
X_4029_ u_bits.i_op2\[17\] u_bits.i_op2\[15\] _1657_ vssd1 vssd1 vccd1 vccd1 _1677_
+ sky130_fd_sc_hd__mux2_1
X_3400_ _0612_ _1174_ vssd1 vssd1 vccd1 vccd1 o_add[16] sky130_fd_sc_hd__xnor2_4
X_4380_ u_bits.i_op2\[11\] _1892_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__xnor2_1
X_3331_ _0731_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__buf_2
X_3262_ _0697_ u_bits.i_op2\[29\] vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__nand2_1
X_5001_ _2056_ _2348_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__or2b_1
X_3193_ u_muldiv.dividend\[27\] _0742_ _0743_ u_muldiv.o_div\[27\] _0744_ vssd1 vssd1
+ vccd1 vccd1 _0994_ sky130_fd_sc_hd__a221o_1
X_5765_ clknet_leaf_18_i_clk _0408_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_2977_ _0775_ _0780_ _0784_ _0787_ _0788_ _0789_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__mux4_1
X_5696_ clknet_leaf_29_i_clk _0339_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4716_ u_muldiv.divisor\[39\] u_muldiv.divisor\[38\] u_muldiv.divisor\[37\] u_muldiv.divisor\[36\]
+ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__or4_1
X_4647_ u_muldiv.divisor\[5\] u_muldiv.dividend\[5\] vssd1 vssd1 vccd1 vccd1 _2070_
+ sky130_fd_sc_hd__and2b_1
X_4578_ _2013_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__clkbuf_1
X_3529_ _0916_ _0788_ _0917_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__or3b_1
X_2900_ _0629_ _0631_ _0686_ _0713_ _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__a221o_1
X_3880_ _1588_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__clkbuf_1
X_2831_ u_bits.i_op1\[19\] vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__buf_4
X_5550_ clknet_leaf_8_i_clk _0197_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_2762_ _0515_ _0520_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__or2b_2
X_4501_ u_muldiv.mul\[10\] u_muldiv.mul\[11\] _1978_ vssd1 vssd1 vccd1 vccd1 _1982_
+ sky130_fd_sc_hd__mux2_1
X_5481_ clknet_leaf_38_i_clk _0129_ vssd1 vssd1 vccd1 vccd1 u_mux.i_add_override sky130_fd_sc_hd__dfxtp_1
X_2693_ _0500_ _0501_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__and2_1
X_4432_ u_bits.i_op2\[21\] u_bits.i_op2\[20\] _1927_ vssd1 vssd1 vccd1 vccd1 _1934_
+ sky130_fd_sc_hd__or3_1
X_4363_ _1406_ _1873_ _1846_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__o21ai_1
X_3314_ u_muldiv.dividend\[31\] _0721_ _0723_ u_muldiv.o_div\[31\] _0724_ vssd1 vssd1
+ vccd1 vccd1 _1107_ sky130_fd_sc_hd__a221o_1
X_4294_ csr_data\[29\] i_csr_data[29] _1595_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__mux2_1
X_3245_ _0458_ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__xnor2_1
X_3176_ _0617_ _0638_ _0978_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__and3_1
X_5748_ clknet_leaf_24_i_clk _0391_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_5679_ clknet_leaf_31_i_clk _0322_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[25\] sky130_fd_sc_hd__dfxtp_1
X_3030_ _0838_ _0840_ _0760_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__mux2_1
X_4981_ _2070_ _2057_ _2069_ _1826_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__o31ai_1
X_3932_ _0646_ i_op1[19] _1610_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__mux2_1
X_3863_ o_add[21] _1579_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__and2_1
X_5602_ clknet_leaf_32_i_clk _0249_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[19\] sky130_fd_sc_hd__dfxtp_1
X_2814_ _0628_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__buf_2
X_5533_ clknet_leaf_14_i_clk _0181_ vssd1 vssd1 vccd1 vccd1 csr_data\[17\] sky130_fd_sc_hd__dfxtp_1
X_3794_ u_bits.i_op2\[15\] _0654_ _0637_ _1515_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__o22a_1
X_2745_ u_bits.i_op1\[6\] u_muldiv.add_prev\[6\] _0448_ vssd1 vssd1 vccd1 vccd1 _0560_
+ sky130_fd_sc_hd__mux2_2
X_5464_ clknet_leaf_14_i_clk _0112_ vssd1 vssd1 vccd1 vccd1 o_pc_target[6] sky130_fd_sc_hd__dfxtp_2
X_2676_ u_bits.i_op1\[16\] u_muldiv.add_prev\[16\] _0451_ vssd1 vssd1 vccd1 vccd1
+ _0491_ sky130_fd_sc_hd__mux2_1
X_5395_ clknet_leaf_53_i_clk _0043_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[27\] sky130_fd_sc_hd__dfxtp_4
X_4415_ u_bits.i_op2\[18\] _1920_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__xnor2_1
X_4346_ _1376_ _1863_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__or2_1
X_4277_ _1813_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__clkbuf_1
X_3228_ _0788_ _0705_ _0911_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__o21a_1
X_3159_ _0960_ _0961_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__or2_1
X_4200_ _1773_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__clkbuf_1
X_5180_ _0691_ _2519_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__xnor2_1
X_4131_ _1737_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__clkbuf_1
X_4062_ u_bits.i_op2\[27\] u_bits.i_op2\[25\] _1681_ vssd1 vssd1 vccd1 vccd1 _1700_
+ sky130_fd_sc_hd__mux2_1
X_3013_ _0703_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__inv_2
X_4964_ _2319_ _2320_ _2322_ _2303_ _1827_ vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__o221a_1
X_3915_ _1251_ i_op1[11] _1599_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__mux2_1
X_4895_ _1209_ vssd1 vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__buf_2
X_3846_ _1554_ _1564_ _0446_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__a21o_1
X_3777_ _1499_ _1081_ _0643_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__mux2_1
X_5516_ clknet_leaf_13_i_clk _0164_ vssd1 vssd1 vccd1 vccd1 csr_data\[0\] sky130_fd_sc_hd__dfxtp_1
X_2728_ _0536_ _0537_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__and2_1
X_5447_ clknet_leaf_2_i_clk _0095_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2659_ _0472_ _0473_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__nor2_1
X_5378_ clknet_leaf_47_i_clk _0026_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[10\] sky130_fd_sc_hd__dfxtp_2
X_4329_ _0915_ _1850_ _0923_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__a21oi_1
X_3700_ _1333_ csr_data\[8\] _1388_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__o21ai_1
X_4680_ u_muldiv.dividend\[22\] u_muldiv.divisor\[22\] vssd1 vssd1 vccd1 vccd1 _2103_
+ sky130_fd_sc_hd__and2b_1
X_3631_ _0672_ _1310_ _0637_ _1363_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__o22a_1
X_3562_ _0749_ o_add[1] _1297_ _0747_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__a22o_1
X_5301_ u_muldiv.divisor\[15\] _2614_ _2615_ u_muldiv.divisor\[16\] vssd1 vssd1 vccd1
+ vccd1 _0406_ sky130_fd_sc_hd__a22o_1
X_3493_ o_wdata[4] _1233_ _0799_ u_wr_mux.i_reg_data2\[12\] vssd1 vssd1 vccd1 vccd1
+ _1238_ sky130_fd_sc_hd__a22o_1
X_5232_ _2113_ _2566_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__xor2_1
X_5163_ u_muldiv.dividend\[20\] _2504_ _2485_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__mux2_1
X_4114_ i_res_src[2] _1638_ _1635_ o_res_src[2] vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__a22o_1
X_5094_ _2435_ _2441_ _1877_ vssd1 vssd1 vccd1 vccd1 _2442_ sky130_fd_sc_hd__mux2_1
X_4045_ _1665_ _1686_ _1688_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__a21o_1
X_4947_ _2304_ _2306_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__xnor2_1
X_4878_ u_muldiv.o_div\[29\] _2264_ u_muldiv.o_div\[30\] vssd1 vssd1 vccd1 vccd1 _2272_
+ sky130_fd_sc_hd__o21ai_1
X_3829_ _0628_ _1542_ _1545_ _1548_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_40_i_clk clknet_2_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4801_ u_muldiv.quotient_msk\[14\] u_muldiv.o_div\[14\] _1841_ vssd1 vssd1 vccd1
+ vccd1 _2211_ sky130_fd_sc_hd__o21a_1
X_5781_ clknet_leaf_28_i_clk _0423_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[0\] sky130_fd_sc_hd__dfxtp_1
X_2993_ _0746_ _0805_ _0447_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__a21o_1
X_4732_ u_muldiv.o_div\[1\] _2029_ _2154_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__mux2_1
X_4663_ _2084_ _2085_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__nand2_1
X_3614_ _0670_ _0794_ _0867_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__a21o_1
X_4594_ _1204_ _2019_ _2020_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__nor3_1
X_3545_ _1250_ u_bits.i_op1\[10\] _1251_ _0777_ _0778_ _0783_ vssd1 vssd1 vccd1 vccd1
+ _1281_ sky130_fd_sc_hd__mux4_1
X_3476_ o_wdata[4] u_wr_mux.i_reg_data2\[20\] _1224_ vssd1 vssd1 vccd1 vccd1 _1229_
+ sky130_fd_sc_hd__mux2_1
X_5215_ u_muldiv.dividend\[25\] u_muldiv.dividend\[24\] _2525_ vssd1 vssd1 vccd1 vccd1
+ _2552_ sky130_fd_sc_hd__or3_2
X_5146_ _2084_ _2479_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__nand2_1
X_5077_ _2044_ _2415_ _2425_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__a21oi_1
X_4028_ _1665_ _1674_ _1676_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__a21o_1
X_3330_ _1108_ _1122_ _0446_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__a21o_1
X_5000_ _2355_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__clkbuf_1
X_3261_ _0775_ _1057_ _0784_ _0945_ _0879_ _0789_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__mux4_2
X_3192_ _0993_ vssd1 vssd1 vccd1 vccd1 o_add[27] sky130_fd_sc_hd__inv_2
X_5764_ clknet_leaf_18_i_clk _0407_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_2976_ _0758_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__buf_4
X_5695_ clknet_leaf_29_i_clk _0338_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_4715_ _2136_ u_muldiv.dividend\[30\] _2137_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__a21o_1
X_4646_ _2058_ _2067_ _2068_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__a21boi_1
X_4577_ o_add[25] _2004_ vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__and2_1
X_3528_ _0642_ _0683_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__or2_2
X_3459_ u_wr_mux.i_reg_data2\[12\] o_wdata[4] _0718_ vssd1 vssd1 vccd1 vccd1 _1220_
+ sky130_fd_sc_hd__mux2_1
X_5129_ _1841_ _2466_ _2473_ vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__a21o_1
X_2830_ u_bits.i_op1\[18\] vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__buf_4
X_2761_ _0569_ _0570_ _0562_ _0574_ _0575_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__o221a_2
X_4500_ _1981_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
X_2692_ _0505_ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__nand2_1
X_5480_ clknet_leaf_1_i_clk _0128_ vssd1 vssd1 vccd1 vccd1 u_bits.i_sra sky130_fd_sc_hd__dfxtp_2
X_4431_ u_muldiv.divisor\[52\] _1836_ _1887_ u_muldiv.divisor\[53\] _1933_ vssd1 vssd1
+ vccd1 vccd1 _0218_ sky130_fd_sc_hd__a221o_1
X_4362_ _1877_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__buf_4
X_4293_ _1821_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_1
X_3313_ _0728_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__buf_2
X_3244_ _0461_ u_bits.i_op2\[29\] _0465_ u_bits.i_op1\[29\] vssd1 vssd1 vccd1 vccd1
+ _1042_ sky130_fd_sc_hd__a22o_1
X_3175_ _0689_ u_bits.i_op2\[26\] vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__nand2_1
X_5747_ clknet_leaf_21_i_clk _0390_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[31\]
+ sky130_fd_sc_hd__dfxtp_2
X_2959_ u_bits.i_op1\[21\] _0630_ _0656_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__mux2_1
X_5678_ clknet_leaf_31_i_clk _0321_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[24\] sky130_fd_sc_hd__dfxtp_1
X_4629_ u_muldiv.divisor\[8\] u_muldiv.dividend\[8\] vssd1 vssd1 vccd1 vccd1 _2052_
+ sky130_fd_sc_hd__or2b_1
X_4980_ _2070_ _2057_ _2069_ vssd1 vssd1 vccd1 vccd1 _2337_ sky130_fd_sc_hd__o21a_1
X_3931_ _1617_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__clkbuf_1
X_3862_ _1214_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__clkbuf_2
X_5601_ clknet_leaf_32_i_clk _0248_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[18\] sky130_fd_sc_hd__dfxtp_1
X_2813_ _0627_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__buf_2
X_5532_ clknet_leaf_14_i_clk _0180_ vssd1 vssd1 vccd1 vccd1 csr_data\[16\] sky130_fd_sc_hd__dfxtp_1
X_3793_ u_bits.i_op2\[15\] _0654_ _1267_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__a21oi_1
X_2744_ _0455_ _0558_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__xnor2_4
X_5463_ clknet_leaf_10_i_clk _0111_ vssd1 vssd1 vccd1 vccd1 o_pc_target[5] sky130_fd_sc_hd__dfxtp_2
X_2675_ _0457_ _0489_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__xnor2_1
X_5394_ clknet_leaf_53_i_clk _0042_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[26\] sky130_fd_sc_hd__dfxtp_2
X_4414_ _1850_ _1919_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__nand2_1
X_4345_ _1376_ _1863_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__nand2_1
X_4276_ csr_data\[20\] i_csr_data[20] _1811_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__mux2_1
X_3227_ u_muldiv.mul\[28\] _0740_ _0720_ u_muldiv.mul\[60\] _1025_ vssd1 vssd1 vccd1
+ vccd1 _1026_ sky130_fd_sc_hd__a221o_1
X_3158_ _0960_ _0961_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__nand2_1
X_3089_ _0461_ u_bits.i_op2\[24\] _0465_ u_bits.i_op1\[24\] vssd1 vssd1 vccd1 vccd1
+ _0897_ sky130_fd_sc_hd__a22o_1
X_4130_ o_pc_target[8] i_pc_target[8] _1734_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__mux2_1
X_4061_ _1689_ _1698_ _1699_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__a21o_1
X_3012_ _0779_ _0700_ _0762_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__o21a_1
X_4963_ _0794_ _2321_ vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__xor2_1
X_3914_ _1608_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__clkbuf_1
X_4894_ u_muldiv.quotient_msk\[6\] _1210_ _2279_ u_muldiv.quotient_msk\[7\] vssd1
+ vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__a22o_1
X_3845_ _0749_ o_add[18] _1562_ _1563_ _0453_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__a221o_1
X_3776_ _0818_ _0822_ _1309_ _1314_ _0758_ _0673_ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__mux4_1
X_5515_ clknet_leaf_10_i_clk _0163_ vssd1 vssd1 vccd1 vccd1 o_to_trap sky130_fd_sc_hd__dfxtp_2
X_2727_ _0539_ _0540_ _0541_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__mux2_2
X_5446_ clknet_leaf_9_i_clk _0094_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2658_ u_bits.i_op1\[19\] u_muldiv.add_prev\[19\] _0451_ vssd1 vssd1 vccd1 vccd1
+ _0473_ sky130_fd_sc_hd__mux2_1
X_5377_ clknet_leaf_47_i_clk _0025_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[9\] sky130_fd_sc_hd__dfxtp_2
X_4328_ _1845_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__buf_2
X_4259_ csr_data\[12\] i_csr_data[12] _1800_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__mux2_1
X_3630_ _0687_ _1310_ _1267_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__a21oi_1
X_3561_ _1249_ _1291_ _1296_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__a21bo_1
X_5300_ u_muldiv.divisor\[14\] _2614_ _2615_ u_muldiv.divisor\[15\] vssd1 vssd1 vccd1
+ vccd1 _0405_ sky130_fd_sc_hd__a22o_1
X_3492_ _1192_ u_wr_mux.i_reg_data2\[27\] _1237_ vssd1 vssd1 vccd1 vccd1 o_wdata[27]
+ sky130_fd_sc_hd__a21o_2
X_5231_ _2117_ _2557_ _2114_ vssd1 vssd1 vccd1 vccd1 _2566_ sky130_fd_sc_hd__a21oi_1
X_5162_ _2498_ _2503_ _1877_ vssd1 vssd1 vccd1 vccd1 _2504_ sky130_fd_sc_hd__mux2_1
X_5093_ _2436_ _2438_ _2440_ _2375_ vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__a22o_1
X_4113_ i_res_src[1] _1638_ _1635_ _0730_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__a22o_1
X_4044_ u_bits.i_op2\[20\] _1687_ _1675_ i_op2[20] vssd1 vssd1 vccd1 vccd1 _1688_
+ sky130_fd_sc_hd__a22o_1
X_4946_ _2061_ _2305_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__nand2_1
X_4877_ u_muldiv.o_div\[29\] u_muldiv.o_div\[30\] _2264_ _1207_ vssd1 vssd1 vccd1
+ vccd1 _2271_ sky130_fd_sc_hd__o31a_1
X_3828_ _0672_ _1546_ _1547_ _0800_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__o211a_1
X_3759_ _1333_ csr_data\[12\] _1388_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__o21ai_1
X_5429_ clknet_leaf_1_i_clk _0077_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[20\] sky130_fd_sc_hd__dfxtp_4
X_4800_ u_muldiv.o_div\[13\] u_muldiv.o_div\[14\] _2201_ vssd1 vssd1 vccd1 vccd1 _2210_
+ sky130_fd_sc_hd__or3_2
X_2992_ _0750_ o_add[21] _0802_ _0803_ _0804_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__a221o_1
X_5780_ clknet_leaf_5_i_clk _0003_ vssd1 vssd1 vccd1 vccd1 u_muldiv.add_prev\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_4731_ _2153_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__buf_4
X_4662_ u_muldiv.dividend\[18\] u_muldiv.divisor\[18\] vssd1 vssd1 vccd1 vccd1 _2085_
+ sky130_fd_sc_hd__or2b_1
X_3613_ _0669_ _0788_ _0881_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__or3b_1
X_4593_ op_cnt\[0\] op_cnt\[1\] op_cnt\[2\] vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__and3_1
X_3544_ _0447_ _1279_ _1280_ _1124_ vssd1 vssd1 vccd1 vccd1 o_result[0] sky130_fd_sc_hd__o211a_2
X_3475_ _1228_ vssd1 vssd1 vccd1 vccd1 o_wdata[19] sky130_fd_sc_hd__buf_2
X_5214_ u_muldiv.dividend\[24\] _2525_ u_muldiv.dividend\[25\] vssd1 vssd1 vccd1 vccd1
+ _2551_ sky130_fd_sc_hd__o21ai_1
X_5145_ u_muldiv.dividend\[18\] _2468_ u_muldiv.dividend\[19\] vssd1 vssd1 vccd1 vccd1
+ _2488_ sky130_fd_sc_hd__o21ai_1
X_5076_ _2043_ _2080_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__and2b_1
X_4027_ u_bits.i_op2\[15\] _1663_ _1675_ i_op2[15] vssd1 vssd1 vccd1 vccd1 _1676_
+ sky130_fd_sc_hd__a22o_1
X_4929_ _2062_ _2063_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__nor2_1
X_3260_ _1056_ _1001_ _0774_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__mux2_1
X_3191_ _0991_ _0992_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__xnor2_2
X_5763_ clknet_leaf_19_i_clk _0406_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_4714_ _1834_ u_muldiv.dividend\[31\] vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__and2_1
X_2975_ _0524_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__clkbuf_4
X_5694_ clknet_leaf_27_i_clk _0337_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_4645_ u_muldiv.divisor\[4\] u_muldiv.dividend\[4\] vssd1 vssd1 vccd1 vccd1 _2068_
+ sky130_fd_sc_hd__or2b_1
X_4576_ _0903_ _2007_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__nor2_1
X_3527_ _1249_ _1263_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__nand2_1
X_3458_ _1219_ vssd1 vssd1 vccd1 vccd1 o_wdata[11] sky130_fd_sc_hd__buf_2
X_3389_ _0480_ _1166_ vssd1 vssd1 vccd1 vccd1 o_add[19] sky130_fd_sc_hd__xnor2_4
X_5128_ _1207_ _2467_ _2468_ _2472_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__a31o_1
X_5059_ _1251_ _2409_ vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__xnor2_1
X_2760_ _0554_ _0555_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__nand2_1
X_2691_ u_bits.i_op1\[14\] u_muldiv.add_prev\[14\] _0449_ vssd1 vssd1 vccd1 vccd1
+ _0506_ sky130_fd_sc_hd__mux2_2
X_4430_ _1832_ _1932_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__nor2_1
X_4361_ _1827_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__clkbuf_4
X_4292_ csr_data\[28\] i_csr_data[28] _1811_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__mux2_1
X_3312_ _1104_ _1105_ vssd1 vssd1 vccd1 vccd1 o_add[31] sky130_fd_sc_hd__nor2_4
X_3243_ _0739_ csr_data\[28\] _1041_ _0732_ vssd1 vssd1 vccd1 vccd1 o_result[28] sky130_fd_sc_hd__o211a_2
X_3174_ _0833_ _0976_ _0835_ _0832_ _0879_ _0789_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__mux4_1
X_5746_ clknet_leaf_22_i_clk _0389_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[30\]
+ sky130_fd_sc_hd__dfxtp_4
X_2958_ _0768_ u_bits.i_op2\[21\] _0637_ _0770_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__o22a_1
X_5677_ clknet_leaf_31_i_clk _0320_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[23\] sky130_fd_sc_hd__dfxtp_1
X_4628_ u_muldiv.dividend\[9\] u_muldiv.divisor\[9\] vssd1 vssd1 vccd1 vccd1 _2051_
+ sky130_fd_sc_hd__and2b_1
X_2889_ u_bits.i_op2\[2\] _0703_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__nand2_1
X_4559_ _1157_ _2007_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__nor2_1
X_3930_ _0645_ i_op1[18] _1610_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__mux2_1
X_3861_ _1106_ csr_data\[19\] _1578_ _1124_ vssd1 vssd1 vccd1 vccd1 o_result[19] sky130_fd_sc_hd__o211a_2
X_5600_ clknet_leaf_32_i_clk _0247_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[17\] sky130_fd_sc_hd__dfxtp_1
X_3792_ _0688_ _1512_ _1513_ _1249_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__o211a_1
X_2812_ _0625_ _0626_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__nor2_1
X_5531_ clknet_leaf_14_i_clk _0179_ vssd1 vssd1 vccd1 vccd1 csr_data\[15\] sky130_fd_sc_hd__dfxtp_1
X_2743_ _0448_ u_bits.i_op1\[6\] _0497_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__a31o_1
X_5462_ clknet_leaf_10_i_clk _0110_ vssd1 vssd1 vccd1 vccd1 o_pc_target[4] sky130_fd_sc_hd__dfxtp_2
X_2674_ _0460_ u_bits.i_op2\[16\] u_bits.i_op1\[16\] _0464_ vssd1 vssd1 vccd1 vccd1
+ _0489_ sky130_fd_sc_hd__a22o_1
X_5393_ clknet_leaf_53_i_clk _0041_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[25\] sky130_fd_sc_hd__dfxtp_2
X_4413_ u_bits.i_op2\[16\] u_bits.i_op2\[17\] _1910_ vssd1 vssd1 vccd1 vccd1 _1919_
+ sky130_fd_sc_hd__or3_1
X_4344_ _0688_ _1859_ _1846_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__o21ai_1
X_4275_ _1812_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__clkbuf_1
X_3226_ u_muldiv.dividend\[28\] _0721_ _0723_ u_muldiv.o_div\[28\] _0744_ vssd1 vssd1
+ vccd1 vccd1 _1025_ sky130_fd_sc_hd__a221o_1
X_3157_ u_bits.i_op1\[26\] u_muldiv.add_prev\[26\] _0451_ vssd1 vssd1 vccd1 vccd1
+ _0961_ sky130_fd_sc_hd__mux2_1
X_3088_ _0496_ _0614_ _0736_ _0893_ _0469_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__a2111o_1
X_5729_ clknet_leaf_19_i_clk _0372_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_4060_ u_bits.i_op2\[25\] _1687_ _1596_ i_op2[25] vssd1 vssd1 vccd1 vccd1 _1699_
+ sky130_fd_sc_hd__a22o_1
X_3011_ _0821_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__inv_2
X_4962_ _1255_ _2308_ _2292_ vssd1 vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__o21a_1
X_4893_ u_muldiv.quotient_msk\[5\] _1210_ _2279_ u_muldiv.quotient_msk\[6\] vssd1
+ vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__a22o_1
X_3913_ _1305_ i_op1[10] _1599_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__mux2_1
X_3844_ _0908_ _1556_ _0955_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__a21oi_1
X_3775_ _1497_ _1498_ _0730_ u_pc_sel.i_pc_next\[13\] vssd1 vssd1 vccd1 vccd1 o_result[13]
+ sky130_fd_sc_hd__a2bb2o_2
X_5514_ clknet_leaf_12_i_clk _0162_ vssd1 vssd1 vccd1 vccd1 csr_read sky130_fd_sc_hd__dfxtp_1
X_2726_ _0459_ u_bits.i_op2\[0\] u_bits.i_op1\[0\] _0463_ vssd1 vssd1 vccd1 vccd1
+ _0541_ sky130_fd_sc_hd__a22o_2
X_2657_ _0457_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__xnor2_1
X_5445_ clknet_leaf_2_i_clk _0093_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_5376_ clknet_leaf_47_i_clk _0024_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[8\] sky130_fd_sc_hd__dfxtp_2
X_4327_ u_muldiv.divisor\[32\] _1838_ _1843_ u_muldiv.divisor\[33\] _1849_ vssd1 vssd1
+ vccd1 vccd1 _0198_ sky130_fd_sc_hd__a221o_1
X_4258_ _1803_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__clkbuf_1
X_3209_ _0628_ _1000_ _1009_ _0747_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__o31a_1
X_4189_ u_wr_mux.i_reg_data2\[12\] i_reg_data2[12] _1767_ vssd1 vssd1 vccd1 vccd1
+ _1768_ sky130_fd_sc_hd__mux2_1
X_3560_ _1265_ _1292_ _1295_ _0634_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__o211a_1
X_5230_ u_muldiv.dividend\[26\] _2552_ u_muldiv.dividend\[27\] vssd1 vssd1 vccd1 vccd1
+ _2565_ sky130_fd_sc_hd__o21ai_1
X_3491_ o_wdata[3] _1233_ _0799_ u_wr_mux.i_reg_data2\[11\] vssd1 vssd1 vccd1 vccd1
+ _1237_ sky130_fd_sc_hd__a22o_1
X_5161_ _2500_ _2502_ _2288_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__mux2_1
X_5092_ _0655_ _2439_ vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__xnor2_1
X_4112_ i_res_src[0] _1638_ _1636_ o_res_src[0] vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__a22o_1
X_4043_ _1634_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__buf_2
X_4945_ _2060_ u_muldiv.dividend\[2\] vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__nand2_1
X_4876_ _2167_ _2268_ _2270_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__a21oi_1
X_3827_ _0687_ _1292_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__nand2_1
X_3758_ _1331_ _1479_ _1481_ _1482_ _1357_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__o221a_1
X_2709_ u_bits.i_op2\[3\] vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__buf_4
X_3689_ _1254_ _1262_ _0910_ _0824_ _0670_ _0643_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__mux4_1
X_5428_ clknet_leaf_52_i_clk _0076_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[19\] sky130_fd_sc_hd__dfxtp_4
X_5359_ clknet_leaf_40_i_clk _0007_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[55\] sky130_fd_sc_hd__dfxtp_1
X_2991_ _0452_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__clkbuf_4
X_4730_ u_muldiv.outsign _1206_ _2152_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__a21o_2
X_4661_ u_muldiv.divisor\[18\] u_muldiv.dividend\[18\] vssd1 vssd1 vccd1 vccd1 _2084_
+ sky130_fd_sc_hd__or2b_1
X_3612_ _1342_ _1345_ _0644_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__mux2_1
X_4592_ op_cnt\[0\] op_cnt\[1\] op_cnt\[2\] vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__a21oi_1
X_3543_ _0728_ csr_data\[0\] vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__or2_1
X_3474_ o_wdata[3] u_wr_mux.i_reg_data2\[19\] _1224_ vssd1 vssd1 vccd1 vccd1 _1228_
+ sky130_fd_sc_hd__mux2_1
X_5213_ _2362_ _2548_ _0943_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__a21oi_1
X_5144_ u_muldiv.dividend\[19\] u_muldiv.dividend\[18\] _2468_ vssd1 vssd1 vccd1 vccd1
+ _2487_ sky130_fd_sc_hd__or3_1
X_5075_ u_muldiv.dividend\[12\] _2403_ u_muldiv.dividend\[13\] vssd1 vssd1 vccd1 vccd1
+ _2424_ sky130_fd_sc_hd__o21ai_1
X_4026_ _1595_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__buf_2
X_4928_ _2062_ _2063_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__and2_1
X_4859_ u_muldiv.o_div\[25\] _2250_ u_muldiv.o_div\[26\] vssd1 vssd1 vccd1 vccd1 _2257_
+ sky130_fd_sc_hd__o21ai_1
X_3190_ _0964_ _0967_ _0962_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__a21bo_1
X_5762_ clknet_leaf_19_i_clk _0405_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_2974_ u_bits.i_op1\[9\] _0785_ u_bits.i_op1\[7\] _0786_ _0658_ _0659_ vssd1 vssd1
+ vccd1 vccd1 _0787_ sky130_fd_sc_hd__mux4_2
X_4713_ u_muldiv.divisor\[30\] vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__inv_2
X_5693_ clknet_leaf_27_i_clk _0336_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_4644_ _2059_ _2061_ _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__a31o_1
X_4575_ _0855_ _2007_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__nor2_1
X_3526_ _1254_ _1260_ _0910_ _1262_ _0674_ _0644_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__mux4_1
X_3457_ u_wr_mux.i_reg_data2\[11\] o_wdata[3] _0718_ vssd1 vssd1 vccd1 vccd1 _1219_
+ sky130_fd_sc_hd__mux2_1
X_3388_ _0482_ _1165_ _0478_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__o21a_1
X_5127_ _1880_ _2470_ _2471_ vssd1 vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__and3_1
X_5058_ _1305_ _2394_ _2293_ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__o21a_1
X_4009_ _1634_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__buf_2
X_2690_ _0456_ _0504_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__xnor2_4
X_4360_ u_muldiv.divisor\[38\] _1867_ _1843_ u_muldiv.divisor\[39\] _1876_ vssd1 vssd1
+ vccd1 vccd1 _0204_ sky130_fd_sc_hd__a221o_1
X_3311_ _1070_ _1094_ _1103_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__and3_1
X_4291_ _1820_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
X_3242_ _1026_ _1040_ _0447_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__a21o_1
X_3173_ _0689_ _0943_ _0904_ _0692_ _0651_ _0774_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__mux4_1
X_5745_ clknet_leaf_21_i_clk _0388_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[29\]
+ sky130_fd_sc_hd__dfxtp_2
X_2957_ _0618_ _0639_ _0769_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__and3_1
X_5676_ clknet_leaf_30_i_clk _0319_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[22\] sky130_fd_sc_hd__dfxtp_1
X_2888_ _0702_ u_bits.i_sra vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__nand2_4
X_4627_ _2048_ _2049_ vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__nand2_1
X_4558_ _1214_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__clkbuf_4
X_4489_ _1975_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
X_3509_ _0620_ _1195_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__nand2_1
Xclkbuf_2_3__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3860_ _1567_ _1577_ _0446_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__a21o_1
X_3791_ _0860_ _0911_ _0687_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__a21bo_1
X_2811_ o_funct3[1] o_funct3[0] vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__nand2_2
X_5530_ clknet_leaf_14_i_clk _0178_ vssd1 vssd1 vccd1 vccd1 csr_data\[14\] sky130_fd_sc_hd__dfxtp_1
X_2742_ u_mux.i_group_mux u_bits.i_op2\[6\] vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_53_i_clk clknet_2_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5461_ clknet_leaf_13_i_clk _0109_ vssd1 vssd1 vccd1 vccd1 o_pc_target[3] sky130_fd_sc_hd__dfxtp_2
X_2673_ _0486_ _0487_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__nand2_1
X_4412_ u_muldiv.divisor\[48\] _1867_ _1887_ u_muldiv.divisor\[49\] _1918_ vssd1 vssd1
+ vccd1 vccd1 _0214_ sky130_fd_sc_hd__a221o_1
X_5392_ clknet_leaf_53_i_clk _0040_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[24\] sky130_fd_sc_hd__dfxtp_2
X_4343_ u_muldiv.divisor\[35\] _1838_ _1843_ u_muldiv.divisor\[36\] _1862_ vssd1 vssd1
+ vccd1 vccd1 _0201_ sky130_fd_sc_hd__a221o_1
X_4274_ csr_data\[19\] i_csr_data[19] _1811_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__mux2_1
X_3225_ _1024_ vssd1 vssd1 vccd1 vccd1 o_add[28] sky130_fd_sc_hd__inv_2
X_3156_ _0458_ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__xnor2_1
X_3087_ _0810_ _0852_ _0893_ _0814_ _0894_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__o221a_1
X_5728_ clknet_leaf_20_i_clk _0371_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_3989_ _0688_ _1637_ _1638_ i_op2[4] vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__a22o_1
X_5659_ clknet_leaf_27_i_clk _0302_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[5\] sky130_fd_sc_hd__dfxtp_1
X_3010_ _0648_ _0698_ _0820_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__a21oi_1
X_4961_ _2061_ _2065_ _2318_ _1839_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__a31o_1
X_4892_ u_muldiv.quotient_msk\[4\] _1210_ _2279_ u_muldiv.quotient_msk\[5\] vssd1
+ vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__a22o_1
X_3912_ _1607_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__clkbuf_1
X_3843_ _0858_ _1555_ _1558_ _1561_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__or4_1
X_3774_ _1333_ csr_data\[13\] _1388_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__o21ai_1
X_5513_ clknet_leaf_47_i_clk _0161_ vssd1 vssd1 vccd1 vccd1 u_wr_mux.i_reg_data2\[31\]
+ sky130_fd_sc_hd__dfxtp_2
X_2725_ u_bits.i_op1\[0\] u_muldiv.add_prev\[0\] _0449_ vssd1 vssd1 vccd1 vccd1 _0540_
+ sky130_fd_sc_hd__mux2_2
X_2656_ _0460_ u_bits.i_op2\[19\] u_bits.i_op1\[19\] _0464_ vssd1 vssd1 vccd1 vccd1
+ _0471_ sky130_fd_sc_hd__a22o_1
X_5444_ clknet_leaf_2_i_clk _0092_ vssd1 vssd1 vccd1 vccd1 u_pc_sel.i_pc_next\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_5375_ clknet_leaf_47_i_clk _0023_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[7\] sky130_fd_sc_hd__dfxtp_2
X_4326_ _1832_ _1848_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__nor2_1
X_4257_ csr_data\[11\] i_csr_data[11] _1800_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__mux2_1
X_4188_ _1711_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__clkbuf_4
X_3208_ _0925_ _1003_ _1006_ _0914_ _1008_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__a221o_1
X_3139_ _0943_ _0904_ _0658_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__mux2_1
X_3490_ _1192_ u_wr_mux.i_reg_data2\[26\] _1236_ vssd1 vssd1 vccd1 vccd1 o_wdata[26]
+ sky130_fd_sc_hd__a21o_2
X_5160_ _0630_ _2501_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__xnor2_1
X_5091_ _0776_ _2428_ _2293_ vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__o21ai_1
X_4111_ _1728_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__clkbuf_1
X_4042_ u_bits.i_op2\[21\] u_bits.i_op2\[19\] _1681_ vssd1 vssd1 vccd1 vccd1 _1686_
+ sky130_fd_sc_hd__mux2_1
X_4944_ _2064_ _2289_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__nor2_1
X_4875_ _2161_ _2269_ u_muldiv.o_div\[29\] vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__a21oi_1
X_3826_ _0784_ _0787_ _0780_ _0795_ _0788_ _0789_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__mux4_1
X_3757_ u_muldiv.mul\[12\] _0748_ _1400_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__o21ai_1
X_2708_ _0502_ _0507_ _0510_ _0521_ _0522_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__o221a_1
X_3688_ _1416_ _1417_ _1336_ u_pc_sel.i_pc_next\[7\] vssd1 vssd1 vccd1 vccd1 o_result[7]
+ sky130_fd_sc_hd__a2bb2o_2
X_2639_ _0453_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__buf_2
X_5427_ clknet_leaf_52_i_clk _0075_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op2\[18\] sky130_fd_sc_hd__dfxtp_4
X_5358_ clknet_leaf_40_i_clk _0006_ vssd1 vssd1 vccd1 vccd1 u_muldiv.mul\[54\] sky130_fd_sc_hd__dfxtp_1
X_4309_ _1832_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__clkbuf_4
X_5289_ u_muldiv.divisor\[5\] _2284_ _2285_ u_muldiv.divisor\[6\] vssd1 vssd1 vccd1
+ vccd1 _0396_ sky130_fd_sc_hd__a22o_1
X_2990_ _0629_ _0769_ _0714_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__a21oi_1
X_4660_ _2042_ _2043_ _2081_ _2040_ _2082_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__o311a_1
X_3611_ _0998_ _1344_ _0879_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__mux2_1
X_4591_ op_cnt\[0\] op_cnt\[1\] _2018_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__o21a_1
X_3542_ _1275_ _1276_ _1278_ _0744_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__o2bb2a_1
X_3473_ _1227_ vssd1 vssd1 vccd1 vccd1 o_wdata[18] sky130_fd_sc_hd__buf_2
X_5212_ _0943_ _2362_ _2548_ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__and3_1
X_5143_ _2486_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__clkbuf_1
X_5074_ u_muldiv.dividend\[13\] u_muldiv.dividend\[12\] _2403_ vssd1 vssd1 vccd1 vccd1
+ _2423_ sky130_fd_sc_hd__or3_2
X_4025_ u_bits.i_op2\[16\] u_bits.i_op2\[14\] _1657_ vssd1 vssd1 vccd1 vccd1 _1674_
+ sky130_fd_sc_hd__mux2_1
X_4927_ _1839_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__clkbuf_4
X_4858_ _2181_ _2254_ _2256_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__a21oi_1
X_3809_ u_bits.i_op2\[16\] _0653_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__nand2_1
X_4789_ u_muldiv.o_div\[11\] u_muldiv.o_div\[12\] _2194_ vssd1 vssd1 vccd1 vccd1 _2201_
+ sky130_fd_sc_hd__or3_2
X_5761_ clknet_leaf_19_i_clk _0404_ vssd1 vssd1 vccd1 vccd1 u_muldiv.divisor\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_2973_ u_bits.i_op1\[6\] vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__clkbuf_4
X_4712_ _2030_ _2131_ _2132_ _2133_ _2134_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__a311oi_4
X_5692_ clknet_leaf_26_i_clk _0335_ vssd1 vssd1 vccd1 vccd1 u_muldiv.quotient_msk\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4643_ u_muldiv.divisor\[3\] u_muldiv.dividend\[3\] vssd1 vssd1 vccd1 vccd1 _2066_
+ sky130_fd_sc_hd__and2b_1
X_4574_ _2012_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__clkbuf_1
X_3525_ _1261_ _0693_ _0758_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__mux2_1
X_3456_ _1218_ vssd1 vssd1 vccd1 vccd1 o_wdata[10] sky130_fd_sc_hd__buf_2
X_3387_ _0610_ _1164_ _0494_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__o21a_2
X_5126_ _2385_ _2469_ _0647_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__a21o_1
X_5057_ _2405_ _2406_ _2407_ vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__o21ai_1
X_4008_ u_bits.i_op2\[11\] u_bits.i_op2\[9\] _1657_ vssd1 vssd1 vccd1 vccd1 _1662_
+ sky130_fd_sc_hd__mux2_1
X_3310_ _1070_ _1094_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__a21oi_2
X_4290_ csr_data\[27\] i_csr_data[27] _1811_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__mux2_1
X_3241_ _0750_ o_add[28] _1039_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__a21o_1
X_3172_ _0920_ _0973_ _0974_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__a21o_1
X_5744_ clknet_leaf_21_i_clk _0387_ vssd1 vssd1 vccd1 vccd1 u_muldiv.dividend\[28\]
+ sky130_fd_sc_hd__dfxtp_4
X_2956_ _0768_ u_bits.i_op2\[21\] vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__nand2_1
X_5675_ clknet_leaf_31_i_clk _0318_ vssd1 vssd1 vccd1 vccd1 u_muldiv.o_div\[21\] sky130_fd_sc_hd__dfxtp_1
X_2887_ u_bits.i_op1\[31\] vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__buf_4
X_4626_ u_muldiv.dividend\[10\] u_muldiv.divisor\[10\] vssd1 vssd1 vccd1 vccd1 _2049_
+ sky130_fd_sc_hd__or2b_1
X_4557_ _1150_ _2006_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__nor2_1
X_4488_ u_muldiv.mul\[4\] u_muldiv.mul\[5\] _1584_ vssd1 vssd1 vccd1 vccd1 _1975_
+ sky130_fd_sc_hd__mux2_1
X_3508_ _1244_ _1245_ vssd1 vssd1 vccd1 vccd1 o_wsel[3] sky130_fd_sc_hd__nor2_4
X_3439_ _1206_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__buf_4
X_5109_ u_muldiv.dividend\[15\] _2455_ _2378_ vssd1 vssd1 vccd1 vccd1 _2456_ sky130_fd_sc_hd__mux2_1
X_3790_ _0861_ _0862_ _1339_ _1343_ _0789_ _0674_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__mux4_1
X_2810_ _0617_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__inv_2
X_2741_ _0554_ _0555_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__xnor2_2
X_5460_ clknet_leaf_10_i_clk _0108_ vssd1 vssd1 vccd1 vccd1 o_pc_target[2] sky130_fd_sc_hd__dfxtp_2
X_2672_ u_bits.i_op1\[17\] u_muldiv.add_prev\[17\] _0450_ vssd1 vssd1 vccd1 vccd1
+ _0487_ sky130_fd_sc_hd__mux2_1
X_4411_ _1916_ _1917_ _1833_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__a21oi_1
X_5391_ clknet_leaf_49_i_clk _0039_ vssd1 vssd1 vccd1 vccd1 u_bits.i_op1\[23\] sky130_fd_sc_hd__dfxtp_2
X_4342_ _1860_ _1861_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__nor2_1
X_4273_ _1711_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__clkbuf_4
X_3224_ _1017_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__xnor2_2
.ends

