`timescale 1ps/1ps
module cell_buf
(
    input wire A,
    output wire X
);
    assign X = A;
endmodule
