magic
tech sky130A
magscale 1 2
timestamp 1684271884
<< nwell >>
rect -1115 -145 10 75
<< nmos >>
rect -1005 -595 -975 -500
rect -910 -595 -880 -500
rect -815 -595 -785 -500
rect -720 -595 -690 -500
rect -515 -595 -485 -500
rect -420 -595 -390 -500
rect -325 -595 -295 -500
rect -120 -595 -90 -500
<< pmos >>
rect -1005 -105 -975 35
rect -910 -105 -880 35
rect -815 -105 -785 35
rect -720 -105 -690 35
rect -515 -105 -485 35
rect -420 -105 -390 35
rect -325 -105 -295 35
rect -120 -105 -90 35
<< ndiff >>
rect -1065 -545 -1005 -500
rect -1065 -580 -1055 -545
rect -1020 -580 -1005 -545
rect -1065 -595 -1005 -580
rect -975 -595 -910 -500
rect -880 -595 -815 -500
rect -785 -595 -720 -500
rect -690 -515 -630 -500
rect -690 -550 -675 -515
rect -640 -550 -630 -515
rect -690 -595 -630 -550
rect -575 -545 -515 -500
rect -575 -580 -565 -545
rect -530 -580 -515 -545
rect -575 -595 -515 -580
rect -485 -515 -420 -500
rect -485 -550 -470 -515
rect -435 -550 -420 -515
rect -485 -595 -420 -550
rect -390 -595 -325 -500
rect -295 -515 -235 -500
rect -295 -550 -280 -515
rect -245 -550 -235 -515
rect -295 -595 -235 -550
rect -180 -515 -120 -500
rect -180 -550 -170 -515
rect -135 -550 -120 -515
rect -180 -595 -120 -550
rect -90 -545 -30 -500
rect -90 -580 -75 -545
rect -40 -580 -30 -545
rect -90 -595 -30 -580
<< pdiff >>
rect -1075 20 -1005 35
rect -1075 -15 -1055 20
rect -1020 -15 -1005 20
rect -1075 -105 -1005 -15
rect -975 -55 -910 35
rect -975 -90 -960 -55
rect -925 -90 -910 -55
rect -975 -105 -910 -90
rect -880 20 -815 35
rect -880 -15 -865 20
rect -830 -15 -815 20
rect -880 -105 -815 -15
rect -785 -55 -720 35
rect -785 -90 -770 -55
rect -735 -90 -720 -55
rect -785 -105 -720 -90
rect -690 20 -630 35
rect -690 -15 -675 20
rect -640 -15 -630 20
rect -690 -105 -630 -15
rect -575 -55 -515 35
rect -575 -90 -565 -55
rect -530 -90 -515 -55
rect -575 -105 -515 -90
rect -485 20 -420 35
rect -485 -15 -470 20
rect -435 -15 -420 20
rect -485 -105 -420 -15
rect -390 -55 -325 35
rect -390 -90 -375 -55
rect -340 -90 -325 -55
rect -390 -105 -325 -90
rect -295 20 -235 35
rect -295 -15 -280 20
rect -245 -15 -235 20
rect -295 -105 -235 -15
rect -180 20 -120 35
rect -180 -15 -170 20
rect -135 -15 -120 20
rect -180 -105 -120 -15
rect -90 -105 -30 35
<< ndiffc >>
rect -1055 -580 -1020 -545
rect -675 -550 -640 -515
rect -565 -580 -530 -545
rect -470 -550 -435 -515
rect -280 -550 -245 -515
rect -170 -550 -135 -515
rect -75 -580 -40 -545
<< pdiffc >>
rect -1055 -15 -1020 20
rect -960 -90 -925 -55
rect -865 -15 -830 20
rect -770 -90 -735 -55
rect -675 -15 -640 20
rect -565 -90 -530 -55
rect -470 -15 -435 20
rect -375 -90 -340 -55
rect -280 -15 -245 20
rect -170 -15 -135 20
<< poly >>
rect -1005 35 -975 65
rect -910 35 -880 65
rect -815 35 -785 65
rect -720 35 -690 65
rect -515 35 -485 65
rect -420 35 -390 65
rect -325 35 -295 65
rect -120 35 -90 65
rect -1005 -500 -975 -105
rect -910 -500 -880 -105
rect -815 -500 -785 -105
rect -720 -500 -690 -105
rect -515 -255 -485 -105
rect -540 -285 -485 -255
rect -540 -400 -510 -285
rect -420 -300 -390 -105
rect -325 -205 -295 -105
rect -345 -215 -265 -205
rect -345 -250 -320 -215
rect -285 -250 -265 -215
rect -345 -260 -265 -250
rect -445 -310 -370 -300
rect -445 -345 -425 -310
rect -390 -345 -370 -310
rect -445 -355 -370 -345
rect -540 -410 -465 -400
rect -540 -445 -520 -410
rect -485 -445 -465 -410
rect -540 -455 -465 -445
rect -515 -500 -485 -455
rect -420 -500 -390 -355
rect -325 -400 -295 -260
rect -120 -300 -90 -105
rect -245 -310 -90 -300
rect -245 -345 -225 -310
rect -190 -345 -90 -310
rect -245 -355 -90 -345
rect -325 -410 -170 -400
rect -325 -445 -225 -410
rect -190 -445 -170 -410
rect -325 -455 -170 -445
rect -325 -500 -295 -455
rect -120 -500 -90 -355
rect -1005 -625 -975 -595
rect -910 -625 -880 -595
rect -815 -625 -785 -595
rect -720 -625 -690 -595
rect -515 -630 -485 -595
rect -420 -625 -390 -595
rect -325 -625 -295 -595
rect -120 -625 -90 -595
<< polycont >>
rect -320 -250 -285 -215
rect -425 -345 -390 -310
rect -520 -445 -485 -410
rect -225 -345 -190 -310
rect -225 -445 -190 -410
<< locali >>
rect -1075 20 -10 75
rect -1075 -15 -1055 20
rect -1020 -15 -865 20
rect -830 -15 -675 20
rect -640 0 -470 20
rect -640 -15 -620 0
rect -695 -20 -620 -15
rect -480 -15 -470 0
rect -435 0 -280 20
rect -435 -15 -425 0
rect -575 -55 -520 -35
rect -480 -45 -425 -15
rect -295 -15 -280 0
rect -245 -15 -170 20
rect -135 0 -10 20
rect -135 -15 -120 0
rect -295 -35 -120 -15
rect -980 -90 -960 -55
rect -925 -90 -770 -55
rect -735 -90 -715 -55
rect -980 -110 -715 -90
rect -575 -90 -565 -55
rect -530 -90 -520 -55
rect -575 -205 -520 -90
rect -385 -55 -330 -35
rect -385 -90 -375 -55
rect -340 -90 -330 -55
rect -385 -135 -330 -90
rect -385 -170 -195 -135
rect -575 -215 -265 -205
rect -575 -250 -320 -215
rect -285 -250 -265 -215
rect -575 -260 -265 -250
rect -230 -300 -195 -170
rect -665 -310 -370 -300
rect -665 -345 -425 -310
rect -390 -345 -370 -310
rect -665 -355 -370 -345
rect -315 -310 -170 -300
rect -315 -345 -225 -310
rect -190 -345 -170 -310
rect -315 -355 -170 -345
rect -695 -410 -465 -400
rect -695 -445 -520 -410
rect -485 -445 -465 -410
rect -695 -455 -465 -445
rect -695 -515 -610 -455
rect -315 -495 -280 -355
rect -75 -400 -30 -40
rect -245 -410 -30 -400
rect -245 -445 -225 -410
rect -190 -445 -30 -410
rect -245 -455 -30 -445
rect -1080 -545 -995 -530
rect -1080 -580 -1055 -545
rect -1020 -580 -995 -545
rect -695 -550 -675 -515
rect -640 -550 -610 -515
rect -490 -515 -415 -500
rect -575 -545 -530 -525
rect -1080 -640 -995 -580
rect -575 -580 -565 -545
rect -490 -550 -470 -515
rect -435 -550 -415 -515
rect -490 -570 -415 -550
rect -315 -515 -235 -495
rect -315 -550 -280 -515
rect -245 -550 -235 -515
rect -315 -570 -235 -550
rect -180 -515 -130 -455
rect -180 -550 -170 -515
rect -135 -550 -130 -515
rect -180 -570 -130 -550
rect -75 -545 -30 -525
rect -575 -605 -530 -580
rect -40 -580 -30 -545
rect -75 -605 -30 -580
rect -575 -640 -30 -605
<< viali >>
rect -470 -15 -435 20
rect -280 -15 -245 20
rect -170 -15 -135 20
rect -1055 -580 -1020 -545
rect -470 -550 -435 -515
<< metal1 >>
rect -1075 20 -10 75
rect -1075 -15 -470 20
rect -435 -15 -280 20
rect -245 -15 -170 20
rect -135 -15 -10 20
rect -1075 -65 -10 -15
rect -1065 -515 -10 -500
rect -1065 -530 -470 -515
rect -1080 -545 -470 -530
rect -1080 -580 -1055 -545
rect -1020 -550 -470 -545
rect -435 -550 -10 -515
rect -1020 -580 -10 -550
rect -1080 -640 -10 -580
<< end >>
