
.include ../block_head.spice
.include simulation/rv_fetch.spice

Vi_clk i_clk 0 PULSE 0 {VCC} 0 20ps 20ps 960ps 2000ps

.include simulation/stimuli_rv_fetch.cir

.tran 1p 50n
.print tran format=raw file=simulation/rv_fetch.spice.raw v(*)

.end
