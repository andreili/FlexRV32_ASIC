magic
tech sky130A
magscale 1 2
timestamp 1684582458
<< nwell >>
rect -320 -315 685 -45
rect -320 -1315 685 -1025
<< pwell >>
rect -315 -605 690 -490
rect -1105 -845 -1070 -780
rect -915 -840 -880 -775
rect -725 -840 -690 -775
rect -315 -865 690 -750
<< nmos >>
rect -220 -595 -190 -500
rect -125 -595 -95 -500
rect -30 -595 0 -500
rect 65 -595 95 -500
rect 160 -595 190 -500
rect 255 -595 285 -500
rect 460 -595 490 -500
rect 555 -595 585 -500
rect -1055 -855 -1025 -760
rect -960 -855 -930 -760
rect -865 -855 -835 -760
rect -770 -855 -740 -760
rect -125 -860 -95 -765
rect -30 -860 0 -765
rect 65 -860 95 -765
rect 160 -860 190 -765
rect 255 -860 285 -765
rect 460 -860 490 -765
rect 555 -860 585 -765
<< pmos >>
rect -220 -275 -190 -85
rect -125 -275 -95 -85
rect -30 -275 0 -85
rect 65 -275 95 -85
rect 160 -275 190 -85
rect 255 -275 285 -85
rect 460 -275 490 -85
rect 555 -275 585 -85
rect -125 -1275 -95 -1085
rect -30 -1275 0 -1085
rect 65 -1275 95 -1085
rect 160 -1275 190 -1085
rect 255 -1275 285 -1085
rect 460 -1275 490 -1085
rect 555 -1275 585 -1085
<< ndiff >>
rect -280 -515 -220 -500
rect -280 -580 -270 -515
rect -235 -580 -220 -515
rect -280 -595 -220 -580
rect -190 -595 -125 -500
rect -95 -515 -30 -500
rect -95 -580 -80 -515
rect -45 -580 -30 -515
rect -95 -595 -30 -580
rect 0 -595 65 -500
rect 95 -595 160 -500
rect 190 -595 255 -500
rect 285 -515 345 -500
rect 285 -580 300 -515
rect 335 -580 345 -515
rect 285 -595 345 -580
rect 400 -515 460 -500
rect 400 -580 410 -515
rect 445 -580 460 -515
rect 400 -595 460 -580
rect 490 -595 555 -500
rect 585 -515 645 -500
rect 585 -580 600 -515
rect 635 -580 645 -515
rect 585 -595 645 -580
rect -1120 -780 -1055 -760
rect -1120 -845 -1105 -780
rect -1070 -845 -1055 -780
rect -1120 -855 -1055 -845
rect -1025 -855 -960 -760
rect -930 -775 -865 -760
rect -930 -840 -915 -775
rect -880 -840 -865 -775
rect -930 -855 -865 -840
rect -835 -855 -770 -760
rect -740 -775 -680 -760
rect -740 -840 -725 -775
rect -690 -840 -680 -775
rect -740 -855 -680 -840
rect -185 -780 -125 -765
rect -185 -845 -175 -780
rect -140 -845 -125 -780
rect -185 -860 -125 -845
rect -95 -860 -30 -765
rect 0 -780 65 -765
rect 0 -845 15 -780
rect 50 -845 65 -780
rect 0 -860 65 -845
rect 95 -860 160 -765
rect 190 -860 255 -765
rect 285 -780 345 -765
rect 285 -845 300 -780
rect 335 -845 345 -780
rect 285 -860 345 -845
rect 400 -780 460 -765
rect 400 -845 410 -780
rect 445 -845 460 -780
rect 400 -860 460 -845
rect 490 -860 555 -765
rect 585 -780 645 -765
rect 585 -845 600 -780
rect 635 -845 645 -780
rect 585 -860 645 -845
<< pdiff >>
rect -280 -100 -220 -85
rect -280 -165 -270 -100
rect -235 -165 -220 -100
rect -280 -275 -220 -165
rect -190 -190 -125 -85
rect -190 -255 -175 -190
rect -140 -255 -125 -190
rect -190 -275 -125 -255
rect -95 -100 -30 -85
rect -95 -165 -80 -100
rect -45 -165 -30 -100
rect -95 -275 -30 -165
rect 0 -195 65 -85
rect 0 -260 15 -195
rect 50 -260 65 -195
rect 0 -275 65 -260
rect 95 -100 160 -85
rect 95 -165 110 -100
rect 145 -165 160 -100
rect 95 -275 160 -165
rect 190 -195 255 -85
rect 190 -260 205 -195
rect 240 -260 255 -195
rect 190 -275 255 -260
rect 285 -100 460 -85
rect 285 -165 300 -100
rect 335 -165 410 -100
rect 445 -165 460 -100
rect 285 -275 460 -165
rect 490 -195 555 -85
rect 490 -260 505 -195
rect 540 -260 555 -195
rect 490 -275 555 -260
rect 585 -100 645 -85
rect 585 -165 600 -100
rect 635 -165 645 -100
rect 585 -275 645 -165
rect -185 -1195 -125 -1085
rect -185 -1260 -175 -1195
rect -140 -1260 -125 -1195
rect -185 -1275 -125 -1260
rect -95 -1100 -30 -1085
rect -95 -1165 -80 -1100
rect -45 -1165 -30 -1100
rect -95 -1275 -30 -1165
rect 0 -1195 65 -1085
rect 0 -1260 15 -1195
rect 50 -1260 65 -1195
rect 0 -1275 65 -1260
rect 95 -1100 160 -1085
rect 95 -1165 110 -1100
rect 145 -1165 160 -1100
rect 95 -1275 160 -1165
rect 190 -1195 255 -1085
rect 190 -1260 205 -1195
rect 240 -1260 255 -1195
rect 190 -1275 255 -1260
rect 285 -1100 345 -1085
rect 285 -1165 300 -1100
rect 335 -1165 345 -1100
rect 285 -1275 345 -1165
rect 400 -1195 460 -1085
rect 400 -1260 410 -1195
rect 445 -1260 460 -1195
rect 400 -1275 460 -1260
rect 490 -1100 555 -1085
rect 490 -1165 505 -1100
rect 540 -1165 555 -1100
rect 490 -1275 555 -1165
rect 585 -1195 645 -1085
rect 585 -1260 600 -1195
rect 635 -1260 645 -1195
rect 585 -1275 645 -1260
<< ndiffc >>
rect -270 -580 -235 -515
rect -80 -580 -45 -515
rect 300 -580 335 -515
rect 410 -580 445 -515
rect 600 -580 635 -515
rect -1105 -845 -1070 -780
rect -915 -840 -880 -775
rect -725 -840 -690 -775
rect -175 -845 -140 -780
rect 15 -845 50 -780
rect 300 -845 335 -780
rect 410 -845 445 -780
rect 600 -845 635 -780
<< pdiffc >>
rect -270 -165 -235 -100
rect -175 -255 -140 -190
rect -80 -165 -45 -100
rect 15 -260 50 -195
rect 110 -165 145 -100
rect 205 -260 240 -195
rect 300 -165 335 -100
rect 410 -165 445 -100
rect 505 -260 540 -195
rect 600 -165 635 -100
rect -175 -1260 -140 -1195
rect -80 -1165 -45 -1100
rect 15 -1260 50 -1195
rect 110 -1165 145 -1100
rect 205 -1260 240 -1195
rect 300 -1165 335 -1100
rect 410 -1260 445 -1195
rect 505 -1165 540 -1100
rect 600 -1260 635 -1195
<< poly >>
rect -220 -85 -190 -55
rect -125 -85 -95 -55
rect -30 -85 0 -55
rect 65 -85 95 -55
rect 160 -85 190 -55
rect 255 -85 285 -55
rect 460 -85 490 -55
rect 555 -85 585 -55
rect -220 -500 -190 -275
rect -125 -310 -95 -275
rect -140 -330 -85 -310
rect -140 -365 -130 -330
rect -95 -365 -85 -330
rect -140 -385 -85 -365
rect -30 -385 0 -275
rect -125 -500 -95 -385
rect -35 -405 20 -385
rect -35 -440 -25 -405
rect 10 -440 20 -405
rect -35 -460 20 -440
rect -30 -500 0 -460
rect 65 -500 95 -275
rect 160 -385 190 -275
rect 255 -385 285 -275
rect 140 -405 195 -385
rect 140 -440 150 -405
rect 185 -440 195 -405
rect 140 -460 195 -440
rect 240 -405 295 -385
rect 460 -405 490 -275
rect 240 -440 250 -405
rect 285 -440 295 -405
rect 240 -460 295 -440
rect 415 -415 490 -405
rect 415 -450 435 -415
rect 470 -450 490 -415
rect 415 -460 490 -450
rect 160 -500 190 -460
rect 255 -500 285 -460
rect 460 -500 490 -460
rect 555 -500 585 -275
rect -1055 -760 -1025 -520
rect -960 -760 -930 -520
rect -865 -760 -835 -520
rect -770 -760 -740 -520
rect -220 -625 -190 -595
rect -125 -625 -95 -595
rect -30 -625 0 -595
rect -225 -630 -190 -625
rect -230 -635 -190 -630
rect 65 -635 95 -595
rect -285 -655 -190 -635
rect 50 -640 105 -635
rect 40 -645 115 -640
rect -285 -690 -275 -655
rect -240 -660 -195 -655
rect 40 -660 60 -645
rect -240 -665 -200 -660
rect 25 -665 60 -660
rect -240 -670 -205 -665
rect 15 -670 60 -665
rect -240 -675 -210 -670
rect -15 -675 60 -670
rect -240 -680 -215 -675
rect -20 -680 60 -675
rect 95 -680 115 -645
rect -240 -690 -230 -680
rect -285 -710 -230 -690
rect -155 -690 -80 -680
rect -25 -685 115 -680
rect -155 -725 -135 -690
rect -100 -725 -80 -690
rect -155 -735 -80 -725
rect -30 -690 115 -685
rect -30 -695 50 -690
rect -30 -700 35 -695
rect -30 -705 25 -700
rect -30 -710 20 -705
rect -30 -715 10 -710
rect -125 -765 -95 -735
rect -30 -765 0 -715
rect 65 -765 95 -735
rect 160 -765 190 -595
rect 255 -765 285 -595
rect 460 -625 490 -595
rect 555 -635 585 -595
rect 555 -645 630 -635
rect 555 -680 575 -645
rect 610 -680 630 -645
rect 555 -690 630 -680
rect 460 -765 490 -735
rect 555 -765 585 -735
rect -1055 -885 -1025 -855
rect -960 -885 -930 -855
rect -865 -885 -835 -855
rect -770 -885 -740 -855
rect -125 -1085 -95 -860
rect -30 -1085 0 -860
rect 65 -935 95 -860
rect 50 -955 105 -935
rect 50 -990 60 -955
rect 95 -990 105 -955
rect 50 -1010 105 -990
rect 65 -1085 95 -1010
rect 160 -1085 190 -860
rect 255 -1085 285 -860
rect 460 -875 490 -860
rect 395 -905 490 -875
rect 395 -955 450 -905
rect 555 -935 585 -860
rect 395 -990 405 -955
rect 440 -990 450 -955
rect 395 -1040 450 -990
rect 520 -955 585 -935
rect 520 -990 530 -955
rect 565 -990 585 -955
rect 520 -1010 585 -990
rect 395 -1070 490 -1040
rect 460 -1085 490 -1070
rect 555 -1085 585 -1010
rect -125 -1305 -95 -1275
rect -30 -1305 0 -1275
rect 65 -1305 95 -1275
rect 160 -1305 190 -1275
rect 255 -1305 285 -1275
rect 460 -1305 490 -1275
rect 555 -1305 585 -1275
<< polycont >>
rect -130 -365 -95 -330
rect -25 -440 10 -405
rect 150 -440 185 -405
rect 250 -440 285 -405
rect 435 -450 470 -415
rect -275 -690 -240 -655
rect 60 -680 95 -645
rect -135 -725 -100 -690
rect 575 -680 610 -645
rect 60 -990 95 -955
rect 405 -990 440 -955
rect 530 -990 565 -955
<< locali >>
rect -280 -60 645 -45
rect -280 -95 -270 -60
rect -235 -95 15 -60
rect 50 -95 205 -60
rect 240 -95 600 -60
rect 635 -95 645 -60
rect -280 -100 645 -95
rect -280 -165 -270 -100
rect -235 -110 -80 -100
rect -235 -165 -225 -110
rect -280 -185 -225 -165
rect -90 -165 -80 -110
rect -45 -110 110 -100
rect -45 -165 -35 -110
rect -185 -190 -130 -170
rect -90 -185 -35 -165
rect 100 -165 110 -110
rect 145 -110 300 -100
rect 145 -165 155 -110
rect -185 -200 -175 -190
rect -190 -205 -175 -200
rect -195 -210 -175 -205
rect -200 -215 -175 -210
rect -205 -220 -175 -215
rect -210 -255 -175 -220
rect -140 -255 -130 -190
rect -210 -275 -130 -255
rect 5 -195 60 -175
rect 100 -185 155 -165
rect 290 -165 300 -110
rect 335 -165 410 -100
rect 445 -110 600 -100
rect 445 -165 455 -110
rect 5 -260 15 -195
rect 50 -260 60 -195
rect -210 -280 -160 -275
rect -210 -285 -165 -280
rect -210 -290 -170 -285
rect -210 -420 -175 -290
rect 5 -310 60 -260
rect 195 -195 250 -175
rect 290 -185 455 -165
rect 590 -165 600 -110
rect 635 -165 645 -100
rect 195 -260 205 -195
rect 240 -260 250 -195
rect 195 -310 250 -260
rect 495 -195 550 -175
rect 590 -185 645 -165
rect 495 -260 505 -195
rect 540 -260 550 -195
rect 495 -275 550 -260
rect -140 -330 365 -310
rect 495 -315 645 -275
rect -140 -365 -130 -330
rect -95 -350 365 -330
rect -95 -365 -85 -350
rect -140 -385 -85 -365
rect -35 -405 20 -385
rect -35 -420 -25 -405
rect -210 -440 -25 -420
rect 10 -440 20 -405
rect -210 -460 20 -440
rect 140 -405 195 -385
rect 140 -440 150 -405
rect 185 -440 195 -405
rect 140 -460 195 -440
rect 240 -405 295 -385
rect 240 -440 250 -405
rect 285 -440 295 -405
rect 240 -460 295 -440
rect 330 -405 365 -350
rect 530 -405 645 -315
rect 330 -415 490 -405
rect 330 -450 435 -415
rect 470 -450 490 -415
rect 330 -460 490 -450
rect 530 -440 600 -405
rect 635 -440 645 -405
rect -210 -495 -135 -460
rect 330 -495 365 -460
rect 530 -495 645 -440
rect -280 -515 -135 -495
rect -280 -580 -270 -515
rect -235 -580 -135 -515
rect -280 -600 -135 -580
rect -95 -515 230 -495
rect -95 -580 -80 -515
rect -45 -580 230 -515
rect -95 -600 230 -580
rect 285 -515 365 -495
rect 285 -580 300 -515
rect 335 -580 365 -515
rect 285 -600 365 -580
rect 400 -515 450 -495
rect 400 -580 410 -515
rect 445 -580 450 -515
rect -285 -655 -230 -635
rect -285 -690 -275 -655
rect -240 -690 -230 -655
rect -285 -710 -230 -690
rect -170 -680 -135 -600
rect -170 -690 -80 -680
rect -170 -725 -135 -690
rect -100 -725 -80 -690
rect -170 -735 -80 -725
rect -1105 -780 -1050 -755
rect -745 -775 -690 -750
rect -1070 -845 -1050 -780
rect -1105 -865 -1050 -845
rect -935 -840 -915 -775
rect -880 -840 -860 -775
rect -935 -885 -860 -840
rect -745 -840 -725 -775
rect -45 -760 5 -600
rect 160 -635 230 -600
rect 400 -635 450 -580
rect 40 -645 120 -640
rect 40 -680 60 -645
rect 95 -680 120 -645
rect 40 -690 120 -680
rect 85 -760 120 -690
rect 160 -725 450 -635
rect -45 -780 50 -760
rect -745 -860 -690 -840
rect -195 -845 -175 -780
rect -140 -845 -120 -780
rect -195 -935 -120 -845
rect -45 -845 15 -780
rect 85 -780 345 -760
rect 85 -810 300 -780
rect -45 -865 50 -845
rect 285 -845 300 -810
rect 335 -845 345 -780
rect 285 -935 345 -845
rect 400 -780 450 -725
rect 400 -845 410 -780
rect 445 -845 450 -780
rect 400 -865 450 -845
rect 485 -515 645 -495
rect 485 -580 600 -515
rect 635 -580 645 -515
rect 485 -600 645 -580
rect 485 -935 520 -600
rect 555 -645 645 -635
rect 555 -680 575 -645
rect 610 -680 645 -645
rect 555 -690 645 -680
rect 600 -775 645 -690
rect 590 -780 645 -775
rect 590 -845 600 -780
rect 635 -845 645 -780
rect 590 -850 645 -845
rect 600 -865 645 -850
rect -195 -955 105 -935
rect -195 -990 60 -955
rect 95 -990 105 -955
rect -195 -1010 105 -990
rect 285 -955 450 -935
rect 285 -990 405 -955
rect 440 -990 450 -955
rect 285 -1010 450 -990
rect 485 -955 575 -935
rect 485 -990 530 -955
rect 565 -990 575 -955
rect 485 -1010 575 -990
rect -95 -1100 -30 -1010
rect 285 -1080 345 -1010
rect 610 -1045 645 -865
rect -95 -1165 -80 -1100
rect -45 -1165 -30 -1100
rect -185 -1195 -130 -1175
rect -95 -1185 -30 -1165
rect 95 -1100 345 -1080
rect 95 -1165 110 -1100
rect 145 -1130 300 -1100
rect 145 -1165 160 -1130
rect -185 -1250 -175 -1195
rect -280 -1260 -175 -1250
rect -140 -1250 -130 -1195
rect 5 -1195 60 -1175
rect 95 -1185 160 -1165
rect 285 -1165 300 -1130
rect 335 -1165 345 -1100
rect 5 -1250 15 -1195
rect -140 -1260 15 -1250
rect 50 -1250 60 -1195
rect 195 -1195 250 -1175
rect 285 -1185 345 -1165
rect 490 -1085 645 -1045
rect 490 -1100 555 -1085
rect 490 -1165 505 -1100
rect 540 -1165 555 -1100
rect 195 -1250 205 -1195
rect 50 -1260 205 -1250
rect 240 -1250 250 -1195
rect 400 -1195 455 -1175
rect 490 -1185 555 -1165
rect 400 -1250 410 -1195
rect 240 -1260 410 -1250
rect 445 -1250 455 -1195
rect 590 -1195 645 -1175
rect 590 -1250 600 -1195
rect 445 -1260 600 -1250
rect 635 -1260 645 -1195
rect -280 -1265 645 -1260
rect -280 -1300 -270 -1265
rect -235 -1300 15 -1265
rect 50 -1300 205 -1265
rect 240 -1300 600 -1265
rect 635 -1300 645 -1265
rect -280 -1315 645 -1300
<< viali >>
rect -270 -95 -235 -60
rect 15 -95 50 -60
rect 205 -95 240 -60
rect 600 -95 635 -60
rect 150 -440 185 -405
rect 250 -440 285 -405
rect 600 -440 635 -405
rect -80 -565 -45 -530
rect 410 -565 445 -530
rect -275 -690 -240 -655
rect 15 -830 50 -795
rect 410 -825 445 -790
rect 600 -830 635 -795
rect -270 -1300 -235 -1265
rect 15 -1300 50 -1265
rect 205 -1300 240 -1265
rect 600 -1300 635 -1265
<< metal1 >>
rect -280 -60 -225 -45
rect -280 -95 -270 -60
rect -235 -95 -225 -60
rect -280 -110 -225 -95
rect 5 -60 60 -45
rect 5 -95 15 -60
rect 50 -95 60 -60
rect 5 -110 60 -95
rect 195 -60 250 -45
rect 195 -95 205 -60
rect 240 -95 250 -60
rect 195 -110 250 -95
rect 590 -60 645 -45
rect 590 -95 600 -60
rect 635 -95 645 -60
rect 590 -110 645 -95
rect 140 -405 195 -385
rect 140 -440 150 -405
rect 185 -440 195 -405
rect 140 -460 195 -440
rect 240 -405 295 -385
rect 240 -440 250 -405
rect 285 -440 295 -405
rect 240 -460 295 -440
rect 590 -405 645 -385
rect 590 -440 600 -405
rect 635 -440 645 -405
rect 590 -460 645 -440
rect -90 -530 -35 -515
rect -90 -565 -80 -530
rect -45 -565 -35 -530
rect -90 -580 -35 -565
rect 400 -530 455 -515
rect 400 -565 410 -530
rect 445 -565 455 -530
rect 400 -580 455 -565
rect -285 -655 -230 -635
rect -285 -690 -275 -655
rect -240 -690 -230 -655
rect -285 -710 -230 -690
rect 5 -795 60 -780
rect 5 -830 15 -795
rect 50 -830 60 -795
rect 5 -845 60 -830
rect 400 -790 455 -775
rect 400 -825 410 -790
rect 445 -825 455 -790
rect 400 -840 455 -825
rect 590 -795 645 -775
rect 590 -830 600 -795
rect 635 -830 645 -795
rect 590 -850 645 -830
rect -280 -1265 -225 -1250
rect -280 -1300 -270 -1265
rect -235 -1300 -225 -1265
rect -280 -1315 -225 -1300
rect 5 -1265 60 -1250
rect 5 -1300 15 -1265
rect 50 -1300 60 -1265
rect 5 -1315 60 -1300
rect 195 -1265 250 -1250
rect 195 -1300 205 -1265
rect 240 -1300 250 -1265
rect 195 -1315 250 -1300
rect 590 -1265 645 -1250
rect 590 -1300 600 -1265
rect 635 -1300 645 -1265
rect 590 -1315 645 -1300
<< labels >>
flabel metal1 -275 -690 -240 -655 5 FreeSans 200 0 0 0 i_data
flabel metal1 600 -440 635 -405 5 FreeSans 200 0 0 0 Qn
flabel metal1 600 -830 635 -795 5 FreeSans 200 0 0 0 Qp
flabel metal1 150 -440 185 -405 5 FreeSans 200 0 0 0 i_clk
flabel metal1 250 -440 285 -405 5 FreeSans 200 0 0 0 i_en
flabel metal1 -270 -95 -235 -60 5 FreeSans 200 0 0 0 VPWR
flabel metal1 -270 -1300 -235 -1265 5 FreeSans 200 0 0 0 VPWR
flabel metal1 -80 -565 -45 -530 5 FreeSans 200 0 0 0 VGND
flabel nwell -270 -1300 -235 -1265 1 FreeSans 200 0 0 0 VPB
flabel nwell -270 -95 -235 -60 1 FreeSans 200 0 0 0 VPB
flabel pwell -80 -565 -45 -530 1 FreeSans 200 0 0 0 VNB
<< end >>
