* NGSPICE file created from rv_decode.ext - technology: sky130A

X_0985_ clknet_3_4__leaf_i_clk _0014_ VSS VSS VCC VCC o_csr_pc_next[15] sky130_fd_sc_hs__dfxtp_2
X_0770_ i_instruction[10] _0283_ _0292_ _0228_ VSS VSS VCC VCC _0293_ sky130_fd_sc_hs__a211o_1
X_0968_ _0455_ VSS VSS VCC VCC _0061_ sky130_fd_sc_hs__clkbuf_1
X_0899_ _0168_ _0403_ _0405_ _0406_ VSS VSS VCC VCC _0407_ sky130_fd_sc_hs__or4_2
X_0822_ _0330_ _0338_ _0174_ VSS VSS VCC VCC _0339_ sky130_fd_sc_hs__a21o_1
X_0753_ i_instruction[3] _0273_ _0277_ i_instruction[8] _0260_ VSS VSS VCC VCC
+ _0278_ sky130_fd_sc_hs__a221o_1
X_0684_ _0214_ VSS VSS VCC VCC _0215_ sky130_fd_sc_hs__buf_4
X_1021_ clknet_3_2__leaf_i_clk _0050_ VSS VSS VCC VCC o_pc[3] sky130_fd_sc_hs__dfxtp_2
X_0805_ _0172_ i_instruction[5] _0213_ _0322_ _0249_ VSS VSS VCC VCC _0323_
+ sky130_fd_sc_hs__a32o_1
X_0736_ i_instruction[12] _0223_ _0236_ _0249_ _0257_ VSS VSS VCC VCC _0262_
+ sky130_fd_sc_hs__a221o_1
X_0667_ _0170_ i_instruction[4] VSS VSS VCC VCC _0198_ sky130_fd_sc_hs__nand2_4
X_0598_ _0146_ VSS VSS VCC VCC _0147_ sky130_fd_sc_hs__buf_8
X_0521_ o_csr_idx[4] VSS VSS VCC VCC _0108_ sky130_fd_sc_hs__inv_2
X_1004_ clknet_3_3__leaf_i_clk _0033_ VSS VSS VCC VCC o_csr_imm[2] sky130_fd_sc_hs__dfxtp_4
X_0719_ _0229_ _0245_ VSS VSS VCC VCC _0246_ sky130_fd_sc_hs__nor2_1
X_0504_ instruction\[5\] _0075_ VSS VSS VCC VCC _0096_ sky130_fd_sc_hs__nand2_1
X_0984_ clknet_3_7__leaf_i_clk _0013_ VSS VSS VCC VCC o_csr_pc_next[14] sky130_fd_sc_hs__dfxtp_2
X_0967_ o_pc[14] i_pc[14] _0446_ VSS VSS VCC VCC _0455_ sky130_fd_sc_hs__mux2_1
X_0898_ _0177_ _0184_ _0196_ _0232_ i_instruction[25] VSS VSS VCC VCC _0406_
+ sky130_fd_sc_hs__a32o_1
X_0821_ _0197_ _0332_ _0336_ _0337_ VSS VSS VCC VCC _0338_ sky130_fd_sc_hs__a211o_1
X_0752_ _0274_ _0276_ VSS VSS VCC VCC _0277_ sky130_fd_sc_hs__nand2_1
X_0683_ _0176_ i_instruction[13] _0169_ VSS VSS VCC VCC _0214_ sky130_fd_sc_hs__and3b_1
X_1020_ clknet_3_0__leaf_i_clk _0049_ VSS VSS VCC VCC o_pc[2] sky130_fd_sc_hs__dfxtp_2
X_0804_ _0192_ _0215_ VSS VSS VCC VCC _0322_ sky130_fd_sc_hs__nor2_1
X_0735_ _0254_ _0260_ _0209_ VSS VSS VCC VCC _0261_ sky130_fd_sc_hs__a21boi_1
X_0666_ _0196_ VSS VSS VCC VCC _0197_ sky130_fd_sc_hs__buf_4
X_0597_ i_stall i_flush VSS VSS VCC VCC _0146_ sky130_fd_sc_hs__nor2_4
X_0520_ _0106_ _0099_ _0107_ VSS VSS VCC VCC o_imm_i[3] sky130_fd_sc_hs__a21oi_4
X_1003_ clknet_3_4__leaf_i_clk _0032_ VSS VSS VCC VCC o_csr_imm[1] sky130_fd_sc_hs__dfxtp_4
X_0718_ i_instruction[1] _0179_ _0224_ _0201_ _0244_ VSS VSS VCC VCC _0245_
+ sky130_fd_sc_hs__o32a_1
X_0649_ _0170_ i_instruction[8] VSS VSS VCC VCC _0182_ sky130_fd_sc_hs__and2_4
X_0503_ _0094_ VSS VSS VCC VCC _0095_ sky130_fd_sc_hs__buf_8
X_0983_ clknet_3_0__leaf_i_clk _0012_ VSS VSS VCC VCC o_csr_pc_next[13] sky130_fd_sc_hs__dfxtp_2
X_0966_ _0454_ VSS VSS VCC VCC _0060_ sky130_fd_sc_hs__clkbuf_1
X_0897_ _0184_ _0194_ _0404_ _0228_ VSS VSS VCC VCC _0405_ sky130_fd_sc_hs__o211a_1
X_0820_ i_instruction[16] _0232_ _0228_ VSS VSS VCC VCC _0337_ sky130_fd_sc_hs__a21o_1
X_0751_ i_instruction[13] _0275_ VSS VSS VCC VCC _0276_ sky130_fd_sc_hs__or2_1
X_0682_ _0211_ _0183_ _0212_ VSS VSS VCC VCC _0213_ sky130_fd_sc_hs__o21a_1
X_0949_ _0445_ VSS VSS VCC VCC _0052_ sky130_fd_sc_hs__clkbuf_1
X_0803_ _0260_ _0302_ VSS VSS VCC VCC _0321_ sky130_fd_sc_hs__or2_4
X_0734_ _0176_ i_instruction[15] i_instruction[13] _0169_ VSS VSS VCC VCC
+ _0260_ sky130_fd_sc_hs__o31ai_4
X_0665_ i_instruction[0] _0180_ VSS VSS VCC VCC _0196_ sky130_fd_sc_hs__nor2_8
X_0596_ _0145_ VSS VSS VCC VCC o_inst_supported sky130_fd_sc_hs__buf_2
X_1002_ clknet_3_3__leaf_i_clk _0031_ VSS VSS VCC VCC o_csr_imm[0] sky130_fd_sc_hs__dfxtp_4
X_0717_ _0179_ _0193_ VSS VSS VCC VCC _0244_ sky130_fd_sc_hs__nand2_1
X_0648_ _0179_ _0180_ VSS VSS VCC VCC _0181_ sky130_fd_sc_hs__nand2_4
X_0579_ o_funct3[1] o_funct3[0] _0132_ VSS VSS VCC VCC _0133_ sky130_fd_sc_hs__and3b_1
X_0502_ _0092_ _0093_ VSS VSS VCC VCC _0094_ sky130_fd_sc_hs__or2_1
X_0982_ clknet_3_7__leaf_i_clk _0011_ VSS VSS VCC VCC o_csr_pc_next[12] sky130_fd_sc_hs__dfxtp_2
X_0965_ o_pc[13] i_pc[13] _0446_ VSS VSS VCC VCC _0454_ sky130_fd_sc_hs__mux2_1
X_0896_ i_instruction[25] _0275_ VSS VSS VCC VCC _0404_ sky130_fd_sc_hs__or2_1
X_0750_ _0176_ _0192_ VSS VSS VCC VCC _0275_ sky130_fd_sc_hs__or2_2
X_0681_ i_instruction[15] i_instruction[13] _0169_ i_instruction[14] VSS VSS VCC
+ VCC _0212_ sky130_fd_sc_hs__and4b_2
X_0948_ o_pc[5] i_pc[5] _0158_ VSS VSS VCC VCC _0445_ sky130_fd_sc_hs__mux2_1
X_0879_ _0172_ i_instruction[5] _0305_ _0388_ _0181_ VSS VSS VCC VCC _0389_
+ sky130_fd_sc_hs__a311o_1
X_0802_ _0165_ o_csr_imm_sel _0319_ _0320_ _0248_ VSS VSS VCC VCC _0030_ sky130_fd_sc_hs__o221a_1
X_0733_ _0187_ _0254_ VSS VSS VCC VCC _0259_ sky130_fd_sc_hs__nand2_1
X_0664_ _0194_ VSS VSS VCC VCC _0195_ sky130_fd_sc_hs__buf_4
X_0595_ o_inst_mret _0144_ VSS VSS VCC VCC _0145_ sky130_fd_sc_hs__or2_1
X_1001_ clknet_3_3__leaf_i_clk _0030_ VSS VSS VCC VCC o_csr_imm_sel sky130_fd_sc_hs__dfxtp_4
X_0716_ _0164_ VSS VSS VCC VCC _0243_ sky130_fd_sc_hs__clkbuf_8
X_0647_ _0171_ i_instruction[1] VSS VSS VCC VCC _0180_ sky130_fd_sc_hs__nand2_8
X_0578_ i_flush _0079_ VSS VSS VCC VCC _0132_ sky130_fd_sc_hs__nor2_8
X_0501_ instruction\[4\] _0068_ instruction\[2\] VSS VSS VCC VCC _0093_ sky130_fd_sc_hs__and3_1
X_0981_ clknet_3_5__leaf_i_clk _0010_ VSS VSS VCC VCC o_csr_pc_next[11] sky130_fd_sc_hs__dfxtp_2
X_0964_ _0453_ VSS VSS VCC VCC _0059_ sky130_fd_sc_hs__clkbuf_1
X_0895_ _0398_ _0401_ _0402_ VSS VSS VCC VCC _0403_ sky130_fd_sc_hs__o21a_1
X_0680_ _0169_ i_instruction[8] VSS VSS VCC VCC _0211_ sky130_fd_sc_hs__nand2_2
X_0947_ _0444_ VSS VSS VCC VCC _0051_ sky130_fd_sc_hs__clkbuf_1
X_0878_ _0177_ i_instruction[23] _0288_ i_instruction[10] _0387_ VSS VSS VCC
+ VCC _0388_ sky130_fd_sc_hs__o221a_1
X_0801_ _0177_ _0233_ _0241_ VSS VSS VCC VCC _0320_ sky130_fd_sc_hs__a21o_1
X_0732_ _0194_ _0255_ _0256_ _0257_ VSS VSS VCC VCC _0258_ sky130_fd_sc_hs__a31o_1
X_0663_ _0193_ VSS VSS VCC VCC _0194_ sky130_fd_sc_hs__buf_4
X_0594_ _0081_ o_csr_read _0141_ _0143_ VSS VSS VCC VCC _0144_ sky130_fd_sc_hs__or4b_4
Xclkbuf_2_3_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_3_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_1000_ clknet_3_4__leaf_i_clk _0029_ VSS VSS VCC VCC o_funct3[1] sky130_fd_sc_hs__dfxtp_4
X_0715_ _0166_ instruction\[5\] _0167_ _0242_ VSS VSS VCC VCC _0021_ sky130_fd_sc_hs__o211a_1
X_0646_ _0170_ i_instruction[0] VSS VSS VCC VCC _0179_ sky130_fd_sc_hs__nand2_4
X_0577_ _0131_ VSS VSS VCC VCC o_alu_ctrl[0] sky130_fd_sc_hs__buf_2
X_0500_ instruction\[3\] _0065_ VSS VSS VCC VCC _0092_ sky130_fd_sc_hs__and2_1
X_0629_ _0163_ VSS VSS VCC VCC _0014_ sky130_fd_sc_hs__clkbuf_1
Xclkbuf_0_i_clk i_clk VSS VSS VCC VCC clknet_0_i_clk sky130_fd_sc_hs__clkbuf_16
X_0980_ clknet_3_7__leaf_i_clk _0009_ VSS VSS VCC VCC o_csr_pc_next[10] sky130_fd_sc_hs__dfxtp_2
X_0963_ o_pc[12] i_pc[12] _0446_ VSS VSS VCC VCC _0453_ sky130_fd_sc_hs__mux2_1
X_0894_ _0184_ _0271_ _0209_ VSS VSS VCC VCC _0402_ sky130_fd_sc_hs__o21a_4
X_0946_ o_pc[4] i_pc[4] _0158_ VSS VSS VCC VCC _0444_ sky130_fd_sc_hs__mux2_1
X_0877_ _0187_ VSS VSS VCC VCC _0387_ sky130_fd_sc_hs__inv_2
X_0800_ _0302_ _0317_ _0318_ _0210_ VSS VSS VCC VCC _0319_ sky130_fd_sc_hs__o31a_1
X_0731_ _0249_ _0221_ _0192_ VSS VSS VCC VCC _0257_ sky130_fd_sc_hs__o21a_1
X_0662_ _0176_ _0192_ VSS VSS VCC VCC _0193_ sky130_fd_sc_hs__nor2_2
X_0593_ _0067_ _0137_ _0142_ _0097_ valid_input VSS VSS VCC VCC _0143_ sky130_fd_sc_hs__o311a_1
X_0929_ _0243_ o_csr_idx[9] _0309_ _0432_ VSS VSS VCC VCC _0045_ sky130_fd_sc_hs__o211a_1
X_0714_ _0230_ _0231_ _0240_ _0241_ VSS VSS VCC VCC _0242_ sky130_fd_sc_hs__a31o_1
X_0645_ _0172_ _0177_ VSS VSS VCC VCC _0178_ sky130_fd_sc_hs__and2_4
X_0576_ o_csr_idx[5] o_csr_imm_sel _0125_ VSS VSS VCC VCC _0131_ sky130_fd_sc_hs__and3_1
X_0628_ o_csr_pc_next[15] i_pc_next[15] _0158_ VSS VSS VCC VCC _0163_ sky130_fd_sc_hs__mux2_1
X_0559_ o_csr_idx[7] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[27] sky130_fd_sc_hs__a21o_2
X_0962_ _0452_ VSS VSS VCC VCC _0058_ sky130_fd_sc_hs__clkbuf_1
X_0893_ _0341_ _0399_ _0400_ VSS VSS VCC VCC _0401_ sky130_fd_sc_hs__or3_2
Xclkbuf_3_2__f_i_clk clknet_2_1_0_i_clk VSS VSS VCC VCC clknet_3_2__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_0945_ _0443_ VSS VSS VCC VCC _0050_ sky130_fd_sc_hs__clkbuf_1
X_0876_ _0210_ _0384_ _0385_ _0228_ VSS VSS VCC VCC _0386_ sky130_fd_sc_hs__a211o_1
X_0730_ _0202_ _0184_ _0201_ VSS VSS VCC VCC _0256_ sky130_fd_sc_hs__a21o_1
X_0661_ _0170_ _0186_ VSS VSS VCC VCC _0192_ sky130_fd_sc_hs__nand2_8
X_0592_ o_csr_imm_sel o_funct3[1] o_funct3[0] _0068_ VSS VSS VCC VCC _0142_
+ sky130_fd_sc_hs__o31a_1
X_0928_ i_instruction[29] _0233_ _0402_ _0429_ _0431_ VSS VSS VCC VCC _0432_
+ sky130_fd_sc_hs__a221o_1
X_0859_ i_instruction[3] _0274_ _0196_ _0370_ _0210_ VSS VSS VCC VCC _0371_
+ sky130_fd_sc_hs__a32o_1
X_0713_ _0168_ VSS VSS VCC VCC _0241_ sky130_fd_sc_hs__buf_4
X_0644_ _0176_ VSS VSS VCC VCC _0177_ sky130_fd_sc_hs__buf_4
X_0575_ o_imm_i[10] _0127_ _0128_ _0130_ o_inst_branch VSS VSS VCC VCC o_alu_ctrl[2]
+ sky130_fd_sc_hs__a311o_4
X_0627_ _0162_ VSS VSS VCC VCC _0013_ sky130_fd_sc_hs__clkbuf_1
X_0558_ o_csr_idx[6] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[26] sky130_fd_sc_hs__a21o_2
X_0489_ _0085_ VSS VSS VCC VCC _0086_ sky130_fd_sc_hs__buf_8
X_0961_ o_pc[11] i_pc[11] _0446_ VSS VSS VCC VCC _0452_ sky130_fd_sc_hs__mux2_1
X_0892_ i_instruction[10] i_instruction[11] _0184_ _0236_ VSS VSS VCC VCC
+ _0400_ sky130_fd_sc_hs__and4b_1
X_0944_ o_pc[3] i_pc[3] _0158_ VSS VSS VCC VCC _0443_ sky130_fd_sc_hs__mux2_1
X_0875_ i_instruction[23] _0232_ _0196_ i_instruction[5] VSS VSS VCC VCC _0385_
+ sky130_fd_sc_hs__a22o_1
X_0660_ _0190_ _0191_ i_flush VSS VSS VCC VCC _0017_ sky130_fd_sc_hs__a21oi_1
X_0591_ _0139_ _0140_ _0137_ VSS VSS VCC VCC _0141_ sky130_fd_sc_hs__a21oi_1
X_0927_ _0228_ _0430_ i_stall VSS VSS VCC VCC _0431_ sky130_fd_sc_hs__a21o_1
X_0858_ _0200_ _0369_ _0341_ VSS VSS VCC VCC _0370_ sky130_fd_sc_hs__o21bai_1
X_0789_ _0134_ VSS VSS VCC VCC _0309_ sky130_fd_sc_hs__buf_4
X_0712_ i_instruction[5] _0233_ _0239_ VSS VSS VCC VCC _0240_ sky130_fd_sc_hs__a21o_1
X_0643_ i_instruction[14] VSS VSS VCC VCC _0176_ sky130_fd_sc_hs__buf_4
X_0574_ o_csr_imm_sel o_funct3[1] _0129_ VSS VSS VCC VCC _0130_ sky130_fd_sc_hs__and3b_1
X_1057_ o_csr_idx[4] VSS VSS VCC VCC o_rs2[4] sky130_fd_sc_hs__buf_2
X_0626_ o_csr_pc_next[14] i_pc_next[14] _0158_ VSS VSS VCC VCC _0162_ sky130_fd_sc_hs__mux2_1
X_0557_ o_csr_idx[5] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[25] sky130_fd_sc_hs__a21o_2
X_0488_ _0064_ instruction\[3\] instruction\[2\] VSS VSS VCC VCC _0085_ sky130_fd_sc_hs__or3b_4
X_0609_ o_csr_pc_next[6] i_pc_next[6] _0147_ VSS VSS VCC VCC _0153_ sky130_fd_sc_hs__mux2_1
X_0960_ _0451_ VSS VSS VCC VCC _0057_ sky130_fd_sc_hs__clkbuf_1
X_0891_ i_instruction[12] _0361_ _0260_ VSS VSS VCC VCC _0399_ sky130_fd_sc_hs__a21o_1
X_0943_ _0442_ VSS VSS VCC VCC _0049_ sky130_fd_sc_hs__clkbuf_1
X_0874_ _0369_ _0383_ _0341_ VSS VSS VCC VCC _0384_ sky130_fd_sc_hs__o21bai_1
X_0590_ _0064_ instruction\[2\] _0074_ VSS VSS VCC VCC _0140_ sky130_fd_sc_hs__a21o_1
X_0926_ _0305_ _0235_ _0194_ i_instruction[29] VSS VSS VCC VCC _0430_ sky130_fd_sc_hs__a22o_1
X_0857_ _0221_ _0361_ VSS VSS VCC VCC _0369_ sky130_fd_sc_hs__nor2_1
X_0788_ _0165_ o_funct3[0] _0307_ _0308_ _0248_ VSS VSS VCC VCC _0028_ sky130_fd_sc_hs__o221a_1
X_0711_ _0186_ _0180_ _0238_ _0179_ VSS VSS VCC VCC _0239_ sky130_fd_sc_hs__o22a_1
X_0642_ _0174_ instruction\[0\] VSS VSS VCC VCC _0175_ sky130_fd_sc_hs__nand2_1
X_0573_ o_csr_idx[5] _0070_ _0128_ VSS VSS VCC VCC _0129_ sky130_fd_sc_hs__o21ai_1
X_1056_ o_csr_idx[3] VSS VSS VCC VCC o_rs2[3] sky130_fd_sc_hs__buf_2
X_0909_ _0243_ o_csr_idx[6] _0309_ _0415_ VSS VSS VCC VCC _0042_ sky130_fd_sc_hs__o211a_1
X_0625_ _0161_ VSS VSS VCC VCC _0012_ sky130_fd_sc_hs__clkbuf_1
X_0556_ o_csr_idx[4] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[24] sky130_fd_sc_hs__a21o_2
X_0487_ _0084_ VSS VSS VCC VCC o_inst_mret sky130_fd_sc_hs__buf_2
X_1039_ o_csr_pc_next[2] VSS VSS VCC VCC o_pc_next[2] sky130_fd_sc_hs__buf_2
X_0608_ _0152_ VSS VSS VCC VCC _0004_ sky130_fd_sc_hs__clkbuf_1
X_0539_ o_csr_idx[11] _0085_ VSS VSS VCC VCC _0118_ sky130_fd_sc_hs__and2_1
X_0890_ _0215_ _0273_ _0333_ i_instruction[2] VSS VSS VCC VCC _0398_ sky130_fd_sc_hs__o31a_1
X_0942_ o_pc[2] i_pc[2] _0158_ VSS VSS VCC VCC _0442_ sky130_fd_sc_hs__mux2_1
X_0873_ _0172_ i_instruction[5] _0237_ VSS VSS VCC VCC _0383_ sky130_fd_sc_hs__a21boi_1
X_0925_ i_instruction[10] _0215_ _0260_ _0428_ VSS VSS VCC VCC _0429_ sky130_fd_sc_hs__a211o_1
X_0856_ _0166_ o_csr_idx[0] _0309_ _0368_ VSS VSS VCC VCC _0036_ sky130_fd_sc_hs__o211a_1
X_0787_ i_instruction[12] _0229_ _0195_ _0168_ VSS VSS VCC VCC _0308_ sky130_fd_sc_hs__a31o_1
X_0710_ _0234_ _0224_ _0237_ i_instruction[1] VSS VSS VCC VCC _0238_ sky130_fd_sc_hs__a31oi_1
X_0641_ _0168_ VSS VSS VCC VCC _0174_ sky130_fd_sc_hs__buf_4
X_0572_ instruction\[2\] _0071_ _0074_ VSS VSS VCC VCC _0128_ sky130_fd_sc_hs__or3_1
X_1055_ o_csr_idx[2] VSS VSS VCC VCC o_rs2[2] sky130_fd_sc_hs__buf_2
X_0908_ _0168_ _0414_ VSS VSS VCC VCC _0415_ sky130_fd_sc_hs__or2_1
X_0839_ _0295_ _0271_ _0321_ _0341_ _0180_ VSS VSS VCC VCC _0353_ sky130_fd_sc_hs__o221a_1
X_0624_ o_csr_pc_next[13] i_pc_next[13] _0158_ VSS VSS VCC VCC _0161_ sky130_fd_sc_hs__mux2_1
X_0555_ o_csr_idx[3] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[23] sky130_fd_sc_hs__a21o_2
X_0486_ o_csr_idx[2] o_csr_idx[1] _0083_ o_csr_idx[9] VSS VSS VCC VCC _0084_
+ sky130_fd_sc_hs__and4b_1
X_1038_ o_csr_pc_next[1] VSS VSS VCC VCC o_pc_next[1] sky130_fd_sc_hs__buf_2
Xclkbuf_3_5__f_i_clk clknet_2_2_0_i_clk VSS VSS VCC VCC clknet_3_5__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_0607_ o_csr_pc_next[5] i_pc_next[5] _0147_ VSS VSS VCC VCC _0152_ sky130_fd_sc_hs__mux2_1
X_0538_ _0092_ _0116_ _0117_ _0086_ VSS VSS VCC VCC o_imm_i[11] sky130_fd_sc_hs__o211a_2
X_0469_ instruction\[3\] instruction\[2\] _0071_ instruction\[6\] VSS VSS VCC
+ VCC _0072_ sky130_fd_sc_hs__or4b_1
X_0941_ _0441_ VSS VSS VCC VCC _0048_ sky130_fd_sc_hs__clkbuf_1
X_0872_ _0174_ _0381_ _0382_ _0248_ VSS VSS VCC VCC _0038_ sky130_fd_sc_hs__o211a_1
X_0924_ i_instruction[12] _0178_ _0400_ VSS VSS VCC VCC _0428_ sky130_fd_sc_hs__a21o_1
X_0855_ _0366_ _0367_ _0174_ VSS VSS VCC VCC _0368_ sky130_fd_sc_hs__a21o_1
X_0786_ _0304_ _0306_ _0289_ VSS VSS VCC VCC _0307_ sky130_fd_sc_hs__o21a_1
X_0640_ _0166_ valid_input _0167_ _0173_ VSS VSS VCC VCC _0015_ sky130_fd_sc_hs__o211a_1
X_0571_ _0086_ _0127_ VSS VSS VCC VCC o_alu_ctrl[4] sky130_fd_sc_hs__nand2_4
X_1054_ o_csr_idx[1] VSS VSS VCC VCC o_rs2[1] sky130_fd_sc_hs__buf_2
X_0907_ _0410_ _0412_ _0413_ _0289_ VSS VSS VCC VCC _0414_ sky130_fd_sc_hs__o22a_1
X_0838_ _0174_ _0347_ _0351_ _0352_ _0134_ VSS VSS VCC VCC _0034_ sky130_fd_sc_hs__o311a_1
X_0769_ _0235_ _0194_ _0291_ _0180_ VSS VSS VCC VCC _0292_ sky130_fd_sc_hs__o211a_1
X_0623_ _0160_ VSS VSS VCC VCC _0011_ sky130_fd_sc_hs__clkbuf_1
X_0554_ o_csr_idx[2] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[22] sky130_fd_sc_hs__a21o_2
X_0485_ _0080_ VSS VSS VCC VCC _0083_ sky130_fd_sc_hs__inv_2
X_1037_ o_csr_read VSS VSS VCC VCC o_inst_csr_req sky130_fd_sc_hs__buf_2
X_0606_ _0151_ VSS VSS VCC VCC _0003_ sky130_fd_sc_hs__clkbuf_1
X_0537_ o_csr_idx[0] _0068_ _0065_ VSS VSS VCC VCC _0117_ sky130_fd_sc_hs__or3b_1
X_0468_ instruction\[5\] _0064_ VSS VSS VCC VCC _0071_ sky130_fd_sc_hs__or2_1
X_0940_ o_pc[1] i_pc[1] _0158_ VSS VSS VCC VCC _0441_ sky130_fd_sc_hs__mux2_1
X_0871_ _0164_ o_csr_idx[2] VSS VSS VCC VCC _0382_ sky130_fd_sc_hs__or2_1
X_0923_ _0243_ o_csr_idx[8] _0309_ _0427_ VSS VSS VCC VCC _0044_ sky130_fd_sc_hs__o211a_1
X_0854_ i_instruction[20] _0195_ _0273_ i_instruction[2] _0289_ VSS VSS VCC
+ VCC _0367_ sky130_fd_sc_hs__a221o_1
X_0785_ i_instruction[12] _0233_ _0197_ _0305_ VSS VSS VCC VCC _0306_ sky130_fd_sc_hs__a22o_1
X_0570_ o_inst_jal _0075_ VSS VSS VCC VCC _0127_ sky130_fd_sc_hs__nor2_4
X_1053_ o_csr_idx[0] VSS VSS VCC VCC o_rs2[0] sky130_fd_sc_hs__buf_2
X_0906_ i_instruction[5] _0221_ _0275_ i_instruction[26] _0259_ VSS VSS VCC
+ VCC _0413_ sky130_fd_sc_hs__o221a_1
X_0837_ _0164_ o_csr_imm[3] VSS VSS VCC VCC _0352_ sky130_fd_sc_hs__or2_1
X_0768_ _0177_ _0270_ VSS VSS VCC VCC _0291_ sky130_fd_sc_hs__or2_1
X_0699_ _0166_ instruction\[4\] _0167_ _0227_ VSS VSS VCC VCC _0020_ sky130_fd_sc_hs__o211a_1
X_0622_ o_csr_pc_next[12] i_pc_next[12] _0158_ VSS VSS VCC VCC _0160_ sky130_fd_sc_hs__mux2_1
X_0553_ o_csr_idx[1] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[21] sky130_fd_sc_hs__a21o_2
X_0484_ _0082_ VSS VSS VCC VCC o_csr_ebreak sky130_fd_sc_hs__buf_2
X_1036_ o_csr_idx[11] VSS VSS VCC VCC o_imm_i[31] sky130_fd_sc_hs__buf_2
X_0605_ o_csr_pc_next[4] i_pc_next[4] _0147_ VSS VSS VCC VCC _0151_ sky130_fd_sc_hs__mux2_1
X_0536_ o_rd[0] o_csr_idx[11] _0097_ VSS VSS VCC VCC _0116_ sky130_fd_sc_hs__mux2_1
X_0467_ instruction\[6\] _0069_ VSS VSS VCC VCC _0070_ sky130_fd_sc_hs__or2_1
X_1019_ clknet_3_5__leaf_i_clk _0048_ VSS VSS VCC VCC o_pc[1] sky130_fd_sc_hs__dfxtp_2
X_0519_ o_rd[3] _0099_ _0086_ VSS VSS VCC VCC _0107_ sky130_fd_sc_hs__o21ai_1
X_0870_ _0289_ _0377_ _0378_ _0380_ VSS VSS VCC VCC _0381_ sky130_fd_sc_hs__o22a_2
X_0999_ clknet_3_3__leaf_i_clk _0028_ VSS VSS VCC VCC o_funct3[0] sky130_fd_sc_hs__dfxtp_4
X_0922_ _0425_ _0426_ _0241_ VSS VSS VCC VCC _0427_ sky130_fd_sc_hs__a21o_1
X_0853_ _0197_ _0359_ _0360_ _0365_ VSS VSS VCC VCC _0366_ sky130_fd_sc_hs__a31o_1
X_0784_ _0187_ VSS VSS VCC VCC _0305_ sky130_fd_sc_hs__buf_4
X_1052_ o_csr_pc_next[15] VSS VSS VCC VCC o_pc_next[15] sky130_fd_sc_hs__buf_2
X_0905_ i_instruction[26] _0207_ _0196_ _0411_ _0206_ VSS VSS VCC VCC _0412_
+ sky130_fd_sc_hs__a221o_1
X_0836_ i_instruction[18] _0233_ _0197_ _0348_ _0350_ VSS VSS VCC VCC _0351_
+ sky130_fd_sc_hs__a221o_1
X_0767_ i_instruction[10] _0288_ _0188_ _0250_ _0289_ VSS VSS VCC VCC _0290_
+ sky130_fd_sc_hs__a2111o_1
X_0698_ _0220_ _0226_ _0174_ VSS VSS VCC VCC _0227_ sky130_fd_sc_hs__a21o_1
X_0621_ _0159_ VSS VSS VCC VCC _0010_ sky130_fd_sc_hs__clkbuf_1
X_0552_ o_csr_idx[0] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[20] sky130_fd_sc_hs__a21o_2
X_0483_ o_csr_idx[0] _0081_ VSS VSS VCC VCC _0082_ sky130_fd_sc_hs__and2_1
X_1035_ o_csr_imm_sel VSS VSS VCC VCC o_funct3[2] sky130_fd_sc_hs__buf_2
X_0819_ _0333_ _0335_ _0272_ VSS VSS VCC VCC _0336_ sky130_fd_sc_hs__o21a_1
X_0604_ _0150_ VSS VSS VCC VCC _0002_ sky130_fd_sc_hs__clkbuf_1
X_0535_ _0115_ VSS VSS VCC VCC o_imm_i[10] sky130_fd_sc_hs__clkbuf_4
X_0466_ instruction\[5\] instruction\[4\] _0063_ VSS VSS VCC VCC _0069_ sky130_fd_sc_hs__nand3_1
X_1018_ clknet_3_6__leaf_i_clk _0047_ VSS VSS VCC VCC o_csr_idx[11] sky130_fd_sc_hs__dfxtp_4
X_0518_ o_csr_idx[3] VSS VSS VCC VCC _0106_ sky130_fd_sc_hs__inv_2
X_0998_ clknet_3_1__leaf_i_clk _0027_ VSS VSS VCC VCC o_rd[4] sky130_fd_sc_hs__dfxtp_2
X_0921_ _0305_ _0284_ _0195_ i_instruction[28] _0289_ VSS VSS VCC VCC _0426_
+ sky130_fd_sc_hs__a221o_1
X_0852_ i_instruction[20] _0232_ _0210_ _0364_ _0206_ VSS VSS VCC VCC _0365_
+ sky130_fd_sc_hs__a221o_1
X_0783_ _0299_ _0300_ _0303_ _0180_ VSS VSS VCC VCC _0304_ sky130_fd_sc_hs__o31a_1
X_1051_ o_csr_pc_next[14] VSS VSS VCC VCC o_pc_next[14] sky130_fd_sc_hs__buf_2
X_0904_ i_instruction[2] _0250_ _0223_ _0249_ VSS VSS VCC VCC _0411_ sky130_fd_sc_hs__a22o_1
X_0835_ _0235_ _0271_ _0349_ _0210_ VSS VSS VCC VCC _0350_ sky130_fd_sc_hs__o211a_1
X_0766_ _0181_ VSS VSS VCC VCC _0289_ sky130_fd_sc_hs__buf_4
X_0697_ _0221_ _0179_ _0222_ _0225_ VSS VSS VCC VCC _0226_ sky130_fd_sc_hs__a31o_1
Xclkbuf_2_2_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_2_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0620_ o_csr_pc_next[11] i_pc_next[11] _0158_ VSS VSS VCC VCC _0159_ sky130_fd_sc_hs__mux2_1
X_0551_ _0118_ VSS VSS VCC VCC _0122_ sky130_fd_sc_hs__buf_8
X_0482_ o_csr_idx[8] _0080_ VSS VSS VCC VCC _0081_ sky130_fd_sc_hs__nor2_2
X_1034_ o_alu_ctrl[3] VSS VSS VCC VCC o_csr_idx[10] sky130_fd_sc_hs__buf_2
X_0818_ i_instruction[8] _0322_ _0334_ _0321_ VSS VSS VCC VCC _0335_ sky130_fd_sc_hs__a211o_1
X_0749_ _0186_ _0221_ VSS VSS VCC VCC _0274_ sky130_fd_sc_hs__or2_2
X_0603_ o_csr_pc_next[3] i_pc_next[3] _0147_ VSS VSS VCC VCC _0150_ sky130_fd_sc_hs__mux2_1
X_0534_ o_alu_ctrl[3] _0085_ VSS VSS VCC VCC _0115_ sky130_fd_sc_hs__and2_1
X_0465_ _0068_ _0067_ VSS VSS VCC VCC o_inst_jal sky130_fd_sc_hs__nor2_4
X_1017_ clknet_3_3__leaf_i_clk _0046_ VSS VSS VCC VCC o_alu_ctrl[3] sky130_fd_sc_hs__dfxtp_4
X_0517_ _0105_ VSS VSS VCC VCC o_imm_i[2] sky130_fd_sc_hs__buf_2
X_0997_ clknet_3_4__leaf_i_clk _0026_ VSS VSS VCC VCC o_rd[3] sky130_fd_sc_hs__dfxtp_2
X_0920_ i_instruction[28] _0233_ _0402_ _0424_ _0228_ VSS VSS VCC VCC _0425_
+ sky130_fd_sc_hs__a221o_1
X_0851_ _0321_ _0341_ _0362_ _0363_ VSS VSS VCC VCC _0364_ sky130_fd_sc_hs__o31a_1
X_0782_ i_instruction[13] _0273_ _0236_ _0301_ _0302_ VSS VSS VCC VCC _0303_
+ sky130_fd_sc_hs__a221o_1
X_1050_ o_csr_pc_next[13] VSS VSS VCC VCC o_pc_next[13] sky130_fd_sc_hs__buf_2
X_0903_ _0401_ _0408_ _0409_ _0402_ VSS VSS VCC VCC _0410_ sky130_fd_sc_hs__o31a_1
X_0834_ _0291_ _0274_ _0302_ _0341_ VSS VSS VCC VCC _0349_ sky130_fd_sc_hs__a211o_1
X_0765_ _0171_ _0186_ VSS VSS VCC VCC _0288_ sky130_fd_sc_hs__and2_1
X_0696_ i_instruction[4] _0207_ _0210_ _0224_ _0206_ VSS VSS VCC VCC _0225_
+ sky130_fd_sc_hs__a221o_1
X_0550_ _0093_ VSS VSS VCC VCC _0121_ sky130_fd_sc_hs__buf_8
X_0481_ o_csr_imm_sel o_funct3[1] o_funct3[0] _0079_ VSS VSS VCC VCC _0080_
+ sky130_fd_sc_hs__or4_1
X_1033_ clknet_3_2__leaf_i_clk _0062_ VSS VSS VCC VCC o_pc[15] sky130_fd_sc_hs__dfxtp_2
X_0817_ _0171_ i_instruction[6] _0212_ VSS VSS VCC VCC _0334_ sky130_fd_sc_hs__and3_1
X_0748_ _0223_ VSS VSS VCC VCC _0273_ sky130_fd_sc_hs__buf_4
X_0679_ _0209_ VSS VSS VCC VCC _0210_ sky130_fd_sc_hs__buf_4
X_0602_ _0149_ VSS VSS VCC VCC _0001_ sky130_fd_sc_hs__clkbuf_1
X_0533_ _0114_ VSS VSS VCC VCC o_imm_i[9] sky130_fd_sc_hs__buf_2
X_0464_ instruction\[3\] VSS VSS VCC VCC _0068_ sky130_fd_sc_hs__clkinv_2
X_1016_ clknet_3_6__leaf_i_clk _0045_ VSS VSS VCC VCC o_csr_idx[9] sky130_fd_sc_hs__dfxtp_4
X_0516_ _0086_ _0104_ VSS VSS VCC VCC _0105_ sky130_fd_sc_hs__and2_1
X_0996_ clknet_3_6__leaf_i_clk _0025_ VSS VSS VCC VCC o_rd[2] sky130_fd_sc_hs__dfxtp_2
X_0850_ _0199_ _0260_ VSS VSS VCC VCC _0363_ sky130_fd_sc_hs__nand2_1
X_0781_ _0176_ i_instruction[13] _0169_ i_instruction[12] VSS VSS VCC VCC
+ _0302_ sky130_fd_sc_hs__and4b_2
X_0979_ clknet_3_7__leaf_i_clk _0008_ VSS VSS VCC VCC o_csr_pc_next[9] sky130_fd_sc_hs__dfxtp_2
X_0902_ _0249_ _0215_ VSS VSS VCC VCC _0409_ sky130_fd_sc_hs__and2_1
X_0833_ _0305_ _0235_ _0325_ i_instruction[10] VSS VSS VCC VCC _0348_ sky130_fd_sc_hs__a22o_1
X_0764_ _0165_ o_rd[2] _0282_ _0287_ _0248_ VSS VSS VCC VCC _0025_ sky130_fd_sc_hs__o221a_1
X_0695_ _0215_ _0223_ VSS VSS VCC VCC _0224_ sky130_fd_sc_hs__nor2_4
X_0480_ instruction\[6\] _0078_ _0076_ VSS VSS VCC VCC _0079_ sky130_fd_sc_hs__nand3_4
X_1032_ clknet_3_5__leaf_i_clk _0061_ VSS VSS VCC VCC o_pc[14] sky130_fd_sc_hs__dfxtp_2
X_0816_ _0211_ _0183_ _0212_ VSS VSS VCC VCC _0333_ sky130_fd_sc_hs__nor3b_4
X_0747_ _0182_ _0271_ _0209_ VSS VSS VCC VCC _0272_ sky130_fd_sc_hs__o21a_1
X_0678_ i_instruction[1] _0179_ VSS VSS VCC VCC _0209_ sky130_fd_sc_hs__nor2_4
X_0601_ o_csr_pc_next[2] i_pc_next[2] _0147_ VSS VSS VCC VCC _0149_ sky130_fd_sc_hs__mux2_1
X_0532_ o_csr_idx[9] _0085_ VSS VSS VCC VCC _0114_ sky130_fd_sc_hs__and2_1
X_0463_ instruction\[3\] _0067_ VSS VSS VCC VCC o_inst_jalr sky130_fd_sc_hs__nor2_4
X_1015_ clknet_3_6__leaf_i_clk _0044_ VSS VSS VCC VCC o_csr_idx[8] sky130_fd_sc_hs__dfxtp_4
X_0515_ o_rd[2] o_csr_idx[2] _0099_ VSS VSS VCC VCC _0104_ sky130_fd_sc_hs__mux2_1
X_0995_ clknet_3_4__leaf_i_clk _0024_ VSS VSS VCC VCC o_rd[1] sky130_fd_sc_hs__dfxtp_2
X_0780_ i_instruction[11] _0235_ VSS VSS VCC VCC _0301_ sky130_fd_sc_hs__nand2_2
X_0978_ clknet_3_0__leaf_i_clk _0007_ VSS VSS VCC VCC o_csr_pc_next[8] sky130_fd_sc_hs__dfxtp_2
X_0901_ _0223_ _0333_ i_instruction[5] VSS VSS VCC VCC _0408_ sky130_fd_sc_hs__o21a_1
X_0832_ i_instruction[18] _0178_ _0315_ VSS VSS VCC VCC _0347_ sky130_fd_sc_hs__o21a_1
X_0763_ i_instruction[9] _0283_ _0285_ _0286_ _0168_ VSS VSS VCC VCC _0287_
+ sky130_fd_sc_hs__a221o_1
X_0694_ _0170_ _0176_ _0186_ VSS VSS VCC VCC _0223_ sky130_fd_sc_hs__and3_4
X_1031_ clknet_3_2__leaf_i_clk _0060_ VSS VSS VCC VCC o_pc[13] sky130_fd_sc_hs__dfxtp_2
X_0815_ _0182_ _0331_ _0178_ VSS VSS VCC VCC _0332_ sky130_fd_sc_hs__a21o_1
X_0746_ _0187_ _0270_ VSS VSS VCC VCC _0271_ sky130_fd_sc_hs__nand2_2
X_0677_ _0206_ _0193_ _0207_ VSS VSS VCC VCC _0208_ sky130_fd_sc_hs__a21o_4
X_0600_ _0148_ VSS VSS VCC VCC _0000_ sky130_fd_sc_hs__clkbuf_1
X_0531_ _0113_ VSS VSS VCC VCC o_imm_i[8] sky130_fd_sc_hs__buf_2
Xclkbuf_3_1__f_i_clk clknet_2_0_0_i_clk VSS VSS VCC VCC clknet_3_1__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_0462_ instruction\[2\] _0065_ VSS VSS VCC VCC _0067_ sky130_fd_sc_hs__nand2_4
X_1014_ clknet_3_4__leaf_i_clk _0043_ VSS VSS VCC VCC o_csr_idx[7] sky130_fd_sc_hs__dfxtp_2
X_0729_ _0254_ _0201_ VSS VSS VCC VCC _0255_ sky130_fd_sc_hs__nand2_1
X_0514_ _0103_ VSS VSS VCC VCC o_imm_i[1] sky130_fd_sc_hs__buf_2
X_0994_ clknet_3_1__leaf_i_clk _0023_ VSS VSS VCC VCC o_rd[0] sky130_fd_sc_hs__dfxtp_4
X_0977_ clknet_3_2__leaf_i_clk _0006_ VSS VSS VCC VCC o_csr_pc_next[7] sky130_fd_sc_hs__dfxtp_2
X_0900_ _0243_ o_csr_idx[5] _0309_ _0407_ VSS VSS VCC VCC _0041_ sky130_fd_sc_hs__o211a_1
X_0831_ _0165_ o_csr_imm[2] _0344_ _0346_ _0248_ VSS VSS VCC VCC _0033_ sky130_fd_sc_hs__o221a_1
X_0762_ i_instruction[4] _0273_ _0277_ i_instruction[9] _0260_ VSS VSS VCC VCC
+ _0286_ sky130_fd_sc_hs__a221o_1
X_0693_ _0192_ _0201_ _0204_ VSS VSS VCC VCC _0222_ sky130_fd_sc_hs__or3_1
X_1030_ clknet_3_5__leaf_i_clk _0059_ VSS VSS VCC VCC o_pc[12] sky130_fd_sc_hs__dfxtp_2
X_0814_ _0192_ _0184_ _0201_ VSS VSS VCC VCC _0331_ sky130_fd_sc_hs__or3b_4
X_0745_ _0171_ i_instruction[13] VSS VSS VCC VCC _0270_ sky130_fd_sc_hs__nand2_1
X_0676_ _0179_ _0180_ VSS VSS VCC VCC _0207_ sky130_fd_sc_hs__nor2_2
X_0530_ o_csr_idx[8] _0085_ VSS VSS VCC VCC _0113_ sky130_fd_sc_hs__and2_1
X_0461_ _0066_ VSS VSS VCC VCC o_inst_branch sky130_fd_sc_hs__clkbuf_4
X_1013_ clknet_3_6__leaf_i_clk _0042_ VSS VSS VCC VCC o_csr_idx[6] sky130_fd_sc_hs__dfxtp_4
X_0728_ _0171_ _0249_ VSS VSS VCC VCC _0254_ sky130_fd_sc_hs__nand2_1
X_0659_ _0174_ instruction\[1\] VSS VSS VCC VCC _0191_ sky130_fd_sc_hs__nand2_1
X_0513_ _0086_ _0102_ VSS VSS VCC VCC _0103_ sky130_fd_sc_hs__and2_1
X_0993_ clknet_3_1__leaf_i_clk _0022_ VSS VSS VCC VCC instruction\[6\] sky130_fd_sc_hs__dfxtp_4
X_0976_ clknet_3_0__leaf_i_clk _0005_ VSS VSS VCC VCC o_csr_pc_next[6] sky130_fd_sc_hs__dfxtp_2
X_0830_ _0229_ _0345_ _0241_ VSS VSS VCC VCC _0346_ sky130_fd_sc_hs__a21o_1
X_0761_ _0284_ _0271_ _0209_ VSS VSS VCC VCC _0285_ sky130_fd_sc_hs__o21a_1
X_0692_ _0170_ _0176_ VSS VSS VCC VCC _0221_ sky130_fd_sc_hs__nand2_8
X_0959_ o_pc[10] i_pc[10] _0446_ VSS VSS VCC VCC _0451_ sky130_fd_sc_hs__mux2_1
X_0813_ _0177_ _0182_ _0195_ i_instruction[16] _0189_ VSS VSS VCC VCC _0330_
+ sky130_fd_sc_hs__a221o_1
X_0744_ i_instruction[8] _0194_ _0250_ i_instruction[3] _0268_ VSS VSS VCC VCC
+ _0269_ sky130_fd_sc_hs__a221o_1
X_0675_ _0179_ _0180_ VSS VSS VCC VCC _0206_ sky130_fd_sc_hs__and2_2
X_0460_ _0063_ _0065_ VSS VSS VCC VCC _0066_ sky130_fd_sc_hs__and2_1
X_1012_ clknet_3_4__leaf_i_clk _0041_ VSS VSS VCC VCC o_csr_idx[5] sky130_fd_sc_hs__dfxtp_4
X_0727_ _0249_ _0194_ _0250_ i_instruction[2] _0252_ VSS VSS VCC VCC _0253_
+ sky130_fd_sc_hs__a221o_1
X_0658_ _0175_ _0190_ i_flush VSS VSS VCC VCC _0016_ sky130_fd_sc_hs__a21oi_1
X_0589_ instruction\[6\] _0138_ instruction\[4\] instruction\[2\] VSS VSS VCC
+ VCC _0139_ sky130_fd_sc_hs__or4b_1
X_0512_ o_rd[1] o_csr_idx[1] _0099_ VSS VSS VCC VCC _0102_ sky130_fd_sc_hs__mux2_4
X_0992_ clknet_3_1__leaf_i_clk _0021_ VSS VSS VCC VCC instruction\[5\] sky130_fd_sc_hs__dfxtp_4
X_0975_ clknet_3_7__leaf_i_clk _0004_ VSS VSS VCC VCC o_csr_pc_next[5] sky130_fd_sc_hs__dfxtp_2
X_0760_ _0172_ i_instruction[9] VSS VSS VCC VCC _0284_ sky130_fd_sc_hs__and2_2
X_0691_ i_instruction[4] _0195_ _0189_ VSS VSS VCC VCC _0220_ sky130_fd_sc_hs__a21o_1
X_0958_ _0450_ VSS VSS VCC VCC _0056_ sky130_fd_sc_hs__clkbuf_1
X_0889_ _0243_ o_csr_idx[4] _0309_ _0397_ VSS VSS VCC VCC _0040_ sky130_fd_sc_hs__o211a_1
X_0812_ _0165_ o_csr_imm[0] _0324_ _0329_ _0248_ VSS VSS VCC VCC _0031_ sky130_fd_sc_hs__o221a_1
X_0743_ _0251_ _0200_ VSS VSS VCC VCC _0268_ sky130_fd_sc_hs__nor2_1
X_0674_ _0201_ _0204_ VSS VSS VCC VCC _0205_ sky130_fd_sc_hs__nor2_1
X_1011_ clknet_3_4__leaf_i_clk _0040_ VSS VSS VCC VCC o_csr_idx[4] sky130_fd_sc_hs__dfxtp_4
X_0726_ _0251_ _0199_ VSS VSS VCC VCC _0252_ sky130_fd_sc_hs__nor2_1
X_0657_ _0178_ _0189_ _0165_ VSS VSS VCC VCC _0190_ sky130_fd_sc_hs__o21ai_2
X_0588_ o_csr_imm_sel o_funct3[1] instruction\[5\] _0068_ VSS VSS VCC VCC
+ _0138_ sky130_fd_sc_hs__or4_1
X_0511_ _0101_ VSS VSS VCC VCC o_imm_i[0] sky130_fd_sc_hs__buf_2
X_0709_ i_instruction[11] _0235_ _0236_ VSS VSS VCC VCC _0237_ sky130_fd_sc_hs__nand3_2
X_0991_ clknet_3_1__leaf_i_clk _0020_ VSS VSS VCC VCC instruction\[4\] sky130_fd_sc_hs__dfxtp_2
X_0974_ clknet_3_2__leaf_i_clk _0003_ VSS VSS VCC VCC o_csr_pc_next[4] sky130_fd_sc_hs__dfxtp_2
X_0690_ _0166_ instruction\[3\] _0167_ _0219_ VSS VSS VCC VCC _0019_ sky130_fd_sc_hs__o211a_1
Xclkbuf_3_4__f_i_clk clknet_2_2_0_i_clk VSS VSS VCC VCC clknet_3_4__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_0957_ o_pc[9] i_pc[9] _0446_ VSS VSS VCC VCC _0450_ sky130_fd_sc_hs__mux2_1
X_0888_ _0210_ _0393_ _0396_ VSS VSS VCC VCC _0397_ sky130_fd_sc_hs__a21o_1
X_0811_ _0197_ _0259_ _0326_ _0328_ VSS VSS VCC VCC _0329_ sky130_fd_sc_hs__a31o_1
X_0742_ i_instruction[1] _0182_ _0266_ _0168_ VSS VSS VCC VCC _0267_ sky130_fd_sc_hs__a31o_1
X_0673_ _0202_ _0203_ VSS VSS VCC VCC _0204_ sky130_fd_sc_hs__nor2_1
X_1010_ clknet_3_4__leaf_i_clk _0039_ VSS VSS VCC VCC o_csr_idx[3] sky130_fd_sc_hs__dfxtp_4
X_0725_ _0188_ VSS VSS VCC VCC _0251_ sky130_fd_sc_hs__inv_2
X_0656_ _0181_ _0188_ VSS VSS VCC VCC _0189_ sky130_fd_sc_hs__or2_1
X_0587_ instruction\[5\] _0064_ _0063_ _0137_ VSS VSS VCC VCC o_reg_write
+ sky130_fd_sc_hs__a31oi_4
X_0510_ _0095_ _0100_ VSS VSS VCC VCC _0101_ sky130_fd_sc_hs__and2b_2
X_0708_ i_instruction[14] i_instruction[13] i_instruction[15] i_ready VSS VSS
+ VCC VCC _0236_ sky130_fd_sc_hs__and4bb_4
X_0639_ _0168_ _0172_ VSS VSS VCC VCC _0173_ sky130_fd_sc_hs__or2_1
X_0990_ clknet_3_1__leaf_i_clk _0019_ VSS VSS VCC VCC instruction\[3\] sky130_fd_sc_hs__dfxtp_4
X_0973_ clknet_3_0__leaf_i_clk _0002_ VSS VSS VCC VCC o_csr_pc_next[3] sky130_fd_sc_hs__dfxtp_2
X_0956_ _0449_ VSS VSS VCC VCC _0055_ sky130_fd_sc_hs__clkbuf_1
X_0887_ _0172_ _0229_ _0394_ _0395_ VSS VSS VCC VCC _0396_ sky130_fd_sc_hs__a31o_1
X_0810_ _0186_ _0233_ _0327_ i_stall VSS VSS VCC VCC _0328_ sky130_fd_sc_hs__a211o_1
X_0741_ _0221_ _0201_ _0192_ i_instruction[0] VSS VSS VCC VCC _0266_ sky130_fd_sc_hs__a211o_1
X_0672_ _0171_ i_instruction[12] VSS VSS VCC VCC _0203_ sky130_fd_sc_hs__nand2_2
X_0939_ o_csr_idx[11] _0243_ _0439_ _0440_ _0167_ VSS VSS VCC VCC _0047_ sky130_fd_sc_hs__o221a_1
X_0724_ _0186_ _0221_ VSS VSS VCC VCC _0250_ sky130_fd_sc_hs__nor2_2
X_0655_ _0182_ _0183_ _0184_ _0185_ _0187_ VSS VSS VCC VCC _0188_ sky130_fd_sc_hs__o41a_2
X_0586_ instruction\[1\] instruction\[0\] VSS VSS VCC VCC _0137_ sky130_fd_sc_hs__nand2_2
X_0707_ _0171_ i_instruction[10] VSS VSS VCC VCC _0235_ sky130_fd_sc_hs__and2_4
X_0638_ _0171_ VSS VSS VCC VCC _0172_ sky130_fd_sc_hs__buf_4
X_0569_ _0126_ VSS VSS VCC VCC o_alu_ctrl[1] sky130_fd_sc_hs__buf_2
X_0972_ clknet_3_6__leaf_i_clk _0001_ VSS VSS VCC VCC o_csr_pc_next[2] sky130_fd_sc_hs__dfxtp_2
X_0955_ o_pc[8] i_pc[8] _0446_ VSS VSS VCC VCC _0449_ sky130_fd_sc_hs__mux2_1
X_0886_ i_instruction[24] _0232_ _0196_ i_instruction[6] i_stall VSS VSS VCC
+ VCC _0395_ sky130_fd_sc_hs__a221o_1
X_0740_ _0166_ o_rd[0] _0167_ _0265_ VSS VSS VCC VCC _0023_ sky130_fd_sc_hs__o211a_1
X_0671_ _0182_ _0183_ VSS VSS VCC VCC _0202_ sky130_fd_sc_hs__or2_2
X_0938_ i_instruction[31] _0208_ _0241_ VSS VSS VCC VCC _0440_ sky130_fd_sc_hs__a21o_1
X_0869_ _0341_ _0379_ _0210_ VSS VSS VCC VCC _0380_ sky130_fd_sc_hs__o21a_1
Xclkbuf_2_1_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_1_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0723_ i_instruction[7] VSS VSS VCC VCC _0249_ sky130_fd_sc_hs__buf_4
X_0654_ _0176_ _0186_ _0170_ VSS VSS VCC VCC _0187_ sky130_fd_sc_hs__o21ai_4
X_0585_ _0136_ VSS VSS VCC VCC o_csr_clear sky130_fd_sc_hs__buf_2
X_0706_ _0211_ _0183_ _0212_ VSS VSS VCC VCC _0234_ sky130_fd_sc_hs__o21ai_4
X_0637_ _0170_ VSS VSS VCC VCC _0171_ sky130_fd_sc_hs__buf_4
X_0568_ o_csr_idx[5] _0125_ VSS VSS VCC VCC _0126_ sky130_fd_sc_hs__and2_1
X_0499_ _0091_ VSS VSS VCC VCC o_rs1[4] sky130_fd_sc_hs__buf_2
X_0971_ clknet_3_2__leaf_i_clk _0000_ VSS VSS VCC VCC o_csr_pc_next[1] sky130_fd_sc_hs__dfxtp_2
X_0954_ _0448_ VSS VSS VCC VCC _0054_ sky130_fd_sc_hs__clkbuf_1
X_0885_ i_instruction[11] _0192_ _0194_ i_instruction[24] VSS VSS VCC VCC
+ _0394_ sky130_fd_sc_hs__a22o_1
X_0670_ _0185_ _0198_ _0199_ _0200_ VSS VSS VCC VCC _0201_ sky130_fd_sc_hs__nand4b_4
X_0937_ _0321_ _0428_ _0402_ VSS VSS VCC VCC _0439_ sky130_fd_sc_hs__o21a_1
X_0868_ _0198_ _0369_ VSS VSS VCC VCC _0379_ sky130_fd_sc_hs__nor2_1
X_0799_ _0185_ _0301_ _0236_ VSS VSS VCC VCC _0318_ sky130_fd_sc_hs__o21a_1
X_0722_ _0243_ instruction\[6\] _0246_ _0247_ _0248_ VSS VSS VCC VCC _0022_
+ sky130_fd_sc_hs__o221a_1
X_0653_ i_instruction[15] VSS VSS VCC VCC _0186_ sky130_fd_sc_hs__buf_4
X_0584_ o_funct3[1] o_funct3[0] _0132_ VSS VSS VCC VCC _0136_ sky130_fd_sc_hs__and3_1
X_0705_ _0232_ VSS VSS VCC VCC _0233_ sky130_fd_sc_hs__buf_4
X_0636_ _0169_ VSS VSS VCC VCC _0170_ sky130_fd_sc_hs__buf_8
X_0567_ instruction\[6\] _0069_ VSS VSS VCC VCC _0125_ sky130_fd_sc_hs__nor2_1
X_0498_ o_csr_imm[4] _0085_ VSS VSS VCC VCC _0091_ sky130_fd_sc_hs__and2_1
Xclkbuf_3_7__f_i_clk clknet_2_3_0_i_clk VSS VSS VCC VCC clknet_3_7__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_0619_ _0146_ VSS VSS VCC VCC _0158_ sky130_fd_sc_hs__buf_8
X_0970_ _0456_ VSS VSS VCC VCC _0062_ sky130_fd_sc_hs__clkbuf_1
X_0953_ o_pc[7] i_pc[7] _0446_ VSS VSS VCC VCC _0448_ sky130_fd_sc_hs__mux2_1
X_0884_ _0172_ i_instruction[6] _0391_ _0392_ VSS VSS VCC VCC _0393_ sky130_fd_sc_hs__a31o_1
X_0936_ _0165_ o_alu_ctrl[3] _0437_ _0438_ _0167_ VSS VSS VCC VCC _0046_ sky130_fd_sc_hs__o221a_1
X_0867_ i_instruction[22] _0232_ _0197_ i_instruction[4] _0228_ VSS VSS VCC
+ VCC _0378_ sky130_fd_sc_hs__a221o_1
X_0798_ _0234_ _0198_ VSS VSS VCC VCC _0317_ sky130_fd_sc_hs__nor2_1
X_0721_ _0134_ VSS VSS VCC VCC _0248_ sky130_fd_sc_hs__buf_4
X_0652_ i_instruction[5] i_instruction[6] _0169_ VSS VSS VCC VCC _0185_ sky130_fd_sc_hs__o21a_1
X_0583_ _0135_ VSS VSS VCC VCC o_csr_set sky130_fd_sc_hs__buf_2
X_0919_ i_instruction[4] _0333_ _0401_ _0423_ VSS VSS VCC VCC _0424_ sky130_fd_sc_hs__a211o_1
X_0704_ _0207_ VSS VSS VCC VCC _0232_ sky130_fd_sc_hs__clkbuf_8
X_0635_ i_ready VSS VSS VCC VCC _0169_ sky130_fd_sc_hs__buf_4
X_0566_ _0092_ _0124_ instruction\[2\] VSS VSS VCC VCC o_op1_src sky130_fd_sc_hs__o21a_2
X_0497_ _0090_ VSS VSS VCC VCC o_rs1[3] sky130_fd_sc_hs__buf_2
X_1049_ o_csr_pc_next[12] VSS VSS VCC VCC o_pc_next[12] sky130_fd_sc_hs__buf_2
X_0618_ _0157_ VSS VSS VCC VCC _0009_ sky130_fd_sc_hs__clkbuf_1
X_0549_ o_csr_imm[4] _0095_ _0120_ VSS VSS VCC VCC o_imm_i[19] sky130_fd_sc_hs__a21o_2
X_0952_ _0447_ VSS VSS VCC VCC _0053_ sky130_fd_sc_hs__clkbuf_1
X_0883_ i_instruction[11] _0215_ _0333_ i_instruction[6] _0341_ VSS VSS VCC
+ VCC _0392_ sky130_fd_sc_hs__a221o_1
X_0935_ i_instruction[30] _0208_ _0241_ VSS VSS VCC VCC _0438_ sky130_fd_sc_hs__a21o_1
X_0866_ i_instruction[22] _0194_ _0273_ i_instruction[4] _0376_ VSS VSS VCC
+ VCC _0377_ sky130_fd_sc_hs__a221o_1
X_0797_ _0166_ o_funct3[1] _0309_ _0316_ VSS VSS VCC VCC _0029_ sky130_fd_sc_hs__o211a_1
X_0720_ i_instruction[6] _0208_ _0241_ VSS VSS VCC VCC _0247_ sky130_fd_sc_hs__a21o_1
X_0651_ _0169_ i_instruction[12] VSS VSS VCC VCC _0184_ sky130_fd_sc_hs__and2_4
X_0582_ o_funct3[0] _0134_ _0123_ o_funct3[1] VSS VSS VCC VCC _0135_ sky130_fd_sc_hs__and4b_1
X_0918_ i_instruction[9] _0215_ _0223_ i_instruction[12] VSS VSS VCC VCC _0423_
+ sky130_fd_sc_hs__a22o_1
X_0849_ _0236_ _0361_ _0199_ VSS VSS VCC VCC _0362_ sky130_fd_sc_hs__o21ba_1
X_0703_ i_instruction[5] _0177_ _0181_ VSS VSS VCC VCC _0231_ sky130_fd_sc_hs__or3_1
X_0634_ i_stall VSS VSS VCC VCC _0168_ sky130_fd_sc_hs__buf_4
X_0565_ _0071_ _0074_ VSS VSS VCC VCC _0124_ sky130_fd_sc_hs__nor2_1
X_0496_ o_csr_imm[3] _0086_ VSS VSS VCC VCC _0090_ sky130_fd_sc_hs__and2_1
X_1048_ o_csr_pc_next[11] VSS VSS VCC VCC o_pc_next[11] sky130_fd_sc_hs__buf_2
X_0617_ o_csr_pc_next[10] i_pc_next[10] _0147_ VSS VSS VCC VCC _0157_ sky130_fd_sc_hs__mux2_1
X_0548_ o_csr_imm[3] _0095_ _0120_ VSS VSS VCC VCC o_imm_i[18] sky130_fd_sc_hs__a21o_2
X_0479_ instruction\[5\] instruction\[4\] _0063_ VSS VSS VCC VCC _0078_ sky130_fd_sc_hs__and3_1
X_0951_ o_pc[6] i_pc[6] _0446_ VSS VSS VCC VCC _0447_ sky130_fd_sc_hs__mux2_1
X_0882_ _0236_ _0301_ _0260_ _0361_ VSS VSS VCC VCC _0391_ sky130_fd_sc_hs__a211o_1
X_0934_ _0435_ _0436_ _0402_ VSS VSS VCC VCC _0437_ sky130_fd_sc_hs__o21a_1
X_0865_ _0186_ _0375_ VSS VSS VCC VCC _0376_ sky130_fd_sc_hs__nor2_1
X_0796_ _0289_ _0314_ _0315_ _0276_ _0168_ VSS VSS VCC VCC _0316_ sky130_fd_sc_hs__a221o_1
X_0650_ i_instruction[7] i_instruction[9] i_instruction[10] i_instruction[11] _0169_
+ VSS VSS VCC VCC _0183_ sky130_fd_sc_hs__o41a_4
X_0581_ i_flush VSS VSS VCC VCC _0134_ sky130_fd_sc_hs__clkinv_2
X_0917_ _0174_ _0421_ _0422_ _0248_ VSS VSS VCC VCC _0043_ sky130_fd_sc_hs__o211a_1
X_0848_ i_instruction[15] i_instruction[13] _0169_ _0176_ VSS VSS VCC VCC
+ _0361_ sky130_fd_sc_hs__and4bb_2
X_0779_ _0172_ i_instruction[5] i_instruction[6] _0236_ VSS VSS VCC VCC _0300_
+ sky130_fd_sc_hs__and4_1
X_0702_ _0229_ _0192_ VSS VSS VCC VCC _0230_ sky130_fd_sc_hs__nand2_1
X_0633_ _0134_ VSS VSS VCC VCC _0167_ sky130_fd_sc_hs__clkbuf_8
X_0564_ o_csr_imm_sel o_funct3[1] o_funct3[0] _0123_ VSS VSS VCC VCC o_csr_read
+ sky130_fd_sc_hs__o31a_4
X_0495_ _0089_ VSS VSS VCC VCC o_rs1[2] sky130_fd_sc_hs__buf_2
X_1047_ o_csr_pc_next[10] VSS VSS VCC VCC o_pc_next[10] sky130_fd_sc_hs__buf_2
X_0616_ _0156_ VSS VSS VCC VCC _0008_ sky130_fd_sc_hs__clkbuf_1
X_0547_ o_csr_imm[2] _0095_ _0120_ VSS VSS VCC VCC o_imm_i[17] sky130_fd_sc_hs__a21o_2
X_0478_ o_res_src[1] o_res_src[2] VSS VSS VCC VCC o_res_src[0] sky130_fd_sc_hs__nor2_4
X_0950_ _0146_ VSS VSS VCC VCC _0446_ sky130_fd_sc_hs__buf_8
X_0881_ _0243_ o_csr_idx[3] _0309_ _0390_ VSS VSS VCC VCC _0039_ sky130_fd_sc_hs__o211a_1
Xclkbuf_3_0__f_i_clk clknet_2_0_0_i_clk VSS VSS VCC VCC clknet_3_0__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_0933_ i_instruction[12] _0178_ _0215_ i_instruction[8] _0260_ VSS VSS VCC
+ VCC _0436_ sky130_fd_sc_hs__a221o_1
X_0864_ _0172_ i_instruction[6] VSS VSS VCC VCC _0375_ sky130_fd_sc_hs__nand2_1
X_0795_ _0181_ _0187_ VSS VSS VCC VCC _0315_ sky130_fd_sc_hs__nor2_2
X_0580_ _0133_ VSS VSS VCC VCC o_csr_write sky130_fd_sc_hs__buf_2
X_0916_ _0164_ o_csr_idx[7] VSS VSS VCC VCC _0422_ sky130_fd_sc_hs__or2_1
X_0847_ _0305_ _0199_ VSS VSS VCC VCC _0360_ sky130_fd_sc_hs__nand2_1
X_0778_ _0234_ _0199_ VSS VSS VCC VCC _0299_ sky130_fd_sc_hs__nor2_1
X_0701_ _0228_ VSS VSS VCC VCC _0229_ sky130_fd_sc_hs__buf_4
X_0632_ _0165_ VSS VSS VCC VCC _0166_ sky130_fd_sc_hs__clkbuf_8
X_0563_ instruction\[6\] _0078_ _0076_ VSS VSS VCC VCC _0123_ sky130_fd_sc_hs__and3_1
X_0494_ o_csr_imm[2] _0086_ VSS VSS VCC VCC _0089_ sky130_fd_sc_hs__and2_1
X_1046_ o_csr_pc_next[9] VSS VSS VCC VCC o_pc_next[9] sky130_fd_sc_hs__buf_2
X_0615_ o_csr_pc_next[9] i_pc_next[9] _0147_ VSS VSS VCC VCC _0156_ sky130_fd_sc_hs__mux2_1
X_0546_ o_csr_imm[1] _0095_ _0120_ VSS VSS VCC VCC o_imm_i[16] sky130_fd_sc_hs__a21o_2
X_0477_ _0067_ VSS VSS VCC VCC o_res_src[1] sky130_fd_sc_hs__clkinv_4
X_1029_ clknet_3_0__leaf_i_clk _0058_ VSS VSS VCC VCC o_pc[11] sky130_fd_sc_hs__dfxtp_2
X_0529_ _0112_ VSS VSS VCC VCC o_imm_i[7] sky130_fd_sc_hs__buf_2
X_0880_ _0386_ _0389_ _0241_ VSS VSS VCC VCC _0390_ sky130_fd_sc_hs__a21o_1
X_0932_ _0235_ _0295_ _0236_ _0434_ VSS VSS VCC VCC _0435_ sky130_fd_sc_hs__o211a_1
X_0863_ _0243_ o_csr_idx[1] _0309_ _0374_ VSS VSS VCC VCC _0037_ sky130_fd_sc_hs__o211a_1
X_0794_ i_instruction[13] _0232_ _0196_ _0177_ _0313_ VSS VSS VCC VCC _0314_
+ sky130_fd_sc_hs__a221o_1
X_0915_ _0417_ _0419_ _0420_ VSS VSS VCC VCC _0421_ sky130_fd_sc_hs__o21a_1
X_0846_ i_instruction[2] _0273_ _0358_ _0193_ _0305_ VSS VSS VCC VCC _0359_
+ sky130_fd_sc_hs__a221o_1
X_0777_ _0174_ _0297_ _0298_ _0248_ VSS VSS VCC VCC _0027_ sky130_fd_sc_hs__o211a_1
X_0700_ _0206_ VSS VSS VCC VCC _0228_ sky130_fd_sc_hs__buf_4
X_0631_ _0164_ VSS VSS VCC VCC _0165_ sky130_fd_sc_hs__buf_4
X_0562_ o_alu_ctrl[3] _0093_ _0118_ VSS VSS VCC VCC o_imm_i[30] sky130_fd_sc_hs__a21o_2
X_0493_ _0088_ VSS VSS VCC VCC o_rs1[1] sky130_fd_sc_hs__buf_2
X_1045_ o_csr_pc_next[8] VSS VSS VCC VCC o_pc_next[8] sky130_fd_sc_hs__buf_2
X_0829_ _0177_ _0284_ _0195_ i_instruction[17] VSS VSS VCC VCC _0345_ sky130_fd_sc_hs__a22o_1
X_0614_ _0155_ VSS VSS VCC VCC _0007_ sky130_fd_sc_hs__clkbuf_1
X_0545_ o_csr_imm[0] _0095_ _0120_ VSS VSS VCC VCC o_imm_i[15] sky130_fd_sc_hs__a21o_2
X_0476_ _0077_ VSS VSS VCC VCC o_res_src[2] sky130_fd_sc_hs__clkbuf_4
X_1028_ clknet_3_5__leaf_i_clk _0057_ VSS VSS VCC VCC o_pc[10] sky130_fd_sc_hs__dfxtp_2
X_0528_ o_csr_idx[7] _0085_ VSS VSS VCC VCC _0112_ sky130_fd_sc_hs__and2_2
X_0459_ instruction\[6\] instruction\[5\] _0064_ VSS VSS VCC VCC _0065_ sky130_fd_sc_hs__and3_1
X_0931_ _0185_ _0301_ _0433_ VSS VSS VCC VCC _0434_ sky130_fd_sc_hs__o21ai_1
X_0862_ _0372_ _0373_ _0241_ VSS VSS VCC VCC _0374_ sky130_fd_sc_hs__a21o_1
X_0793_ _0302_ _0310_ _0312_ _0180_ VSS VSS VCC VCC _0313_ sky130_fd_sc_hs__o31a_1
X_0914_ _0305_ _0182_ _0195_ i_instruction[27] _0181_ VSS VSS VCC VCC _0420_
+ sky130_fd_sc_hs__a221o_1
X_0845_ _0202_ _0203_ _0201_ _0199_ VSS VSS VCC VCC _0358_ sky130_fd_sc_hs__o31ai_1
X_0776_ _0165_ o_rd[4] VSS VSS VCC VCC _0298_ sky130_fd_sc_hs__or2_1
X_0630_ i_stall VSS VSS VCC VCC _0164_ sky130_fd_sc_hs__inv_2
X_0561_ o_csr_idx[9] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[29] sky130_fd_sc_hs__a21o_2
X_0492_ o_csr_imm[1] _0086_ VSS VSS VCC VCC _0088_ sky130_fd_sc_hs__and2_1
X_1044_ o_csr_pc_next[7] VSS VSS VCC VCC o_pc_next[7] sky130_fd_sc_hs__buf_2
X_0828_ i_instruction[17] _0233_ _0197_ _0340_ _0343_ VSS VSS VCC VCC _0344_
+ sky130_fd_sc_hs__a221o_1
X_0759_ _0244_ _0201_ _0180_ VSS VSS VCC VCC _0283_ sky130_fd_sc_hs__o21ba_2
X_0613_ o_csr_pc_next[8] i_pc_next[8] _0147_ VSS VSS VCC VCC _0155_ sky130_fd_sc_hs__mux2_1
X_0544_ o_csr_imm_sel _0095_ _0120_ VSS VSS VCC VCC o_imm_i[14] sky130_fd_sc_hs__a21o_2
X_0475_ instruction\[5\] _0075_ _0076_ VSS VSS VCC VCC _0077_ sky130_fd_sc_hs__and3b_1
X_1027_ clknet_3_7__leaf_i_clk _0056_ VSS VSS VCC VCC o_pc[9] sky130_fd_sc_hs__dfxtp_2
X_0527_ _0111_ VSS VSS VCC VCC o_imm_i[6] sky130_fd_sc_hs__buf_2
X_0458_ instruction\[4\] VSS VSS VCC VCC _0064_ sky130_fd_sc_hs__clkinv_2
X_0930_ i_instruction[10] _0203_ _0295_ VSS VSS VCC VCC _0433_ sky130_fd_sc_hs__o21a_1
X_0861_ i_instruction[21] _0195_ _0273_ i_instruction[3] _0289_ VSS VSS VCC
+ VCC _0373_ sky130_fd_sc_hs__a221o_1
X_0792_ i_instruction[6] _0311_ _0236_ i_instruction[11] VSS VSS VCC VCC _0312_
+ sky130_fd_sc_hs__o211a_1
X_0913_ i_instruction[27] _0232_ _0197_ _0418_ _0228_ VSS VSS VCC VCC _0419_
+ sky130_fd_sc_hs__a221o_1
X_0844_ _0165_ o_csr_imm[4] _0356_ _0357_ _0167_ VSS VSS VCC VCC _0035_ sky130_fd_sc_hs__o221a_1
X_0775_ _0186_ _0289_ _0295_ _0296_ VSS VSS VCC VCC _0297_ sky130_fd_sc_hs__o211a_1
X_0560_ o_csr_idx[8] _0121_ _0122_ VSS VSS VCC VCC o_imm_i[28] sky130_fd_sc_hs__a21o_2
X_0491_ _0087_ VSS VSS VCC VCC o_rs1[0] sky130_fd_sc_hs__buf_2
X_1043_ o_csr_pc_next[6] VSS VSS VCC VCC o_pc_next[6] sky130_fd_sc_hs__buf_2
X_0827_ _0321_ _0341_ _0342_ _0285_ VSS VSS VCC VCC _0343_ sky130_fd_sc_hs__o31a_1
X_0758_ _0280_ _0281_ _0229_ VSS VSS VCC VCC _0282_ sky130_fd_sc_hs__o21a_1
X_0689_ i_instruction[3] _0208_ _0216_ VSS VSS VCC VCC _0219_ sky130_fd_sc_hs__a21o_1
X_0612_ _0154_ VSS VSS VCC VCC _0006_ sky130_fd_sc_hs__clkbuf_1
X_0543_ o_funct3[1] _0095_ _0120_ VSS VSS VCC VCC o_imm_i[13] sky130_fd_sc_hs__a21o_2
X_0474_ instruction\[1\] instruction\[0\] VSS VSS VCC VCC _0076_ sky130_fd_sc_hs__and2_2
X_1026_ clknet_3_0__leaf_i_clk _0055_ VSS VSS VCC VCC o_pc[8] sky130_fd_sc_hs__dfxtp_2
Xclkbuf_3_3__f_i_clk clknet_2_1_0_i_clk VSS VSS VCC VCC clknet_3_3__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_0526_ o_csr_idx[6] _0085_ VSS VSS VCC VCC _0111_ sky130_fd_sc_hs__and2_1
X_0457_ instruction\[3\] instruction\[2\] VSS VSS VCC VCC _0063_ sky130_fd_sc_hs__nor2_2
X_1009_ clknet_3_4__leaf_i_clk _0038_ VSS VSS VCC VCC o_csr_idx[2] sky130_fd_sc_hs__dfxtp_4
X_0509_ o_rd[0] o_inst_store _0099_ o_csr_idx[0] VSS VSS VCC VCC _0100_ sky130_fd_sc_hs__a22o_1
X_0860_ i_instruction[21] _0233_ _0371_ _0229_ VSS VSS VCC VCC _0372_ sky130_fd_sc_hs__a211o_1
X_0791_ _0171_ i_instruction[10] VSS VSS VCC VCC _0311_ sky130_fd_sc_hs__nand2_1
X_0989_ clknet_3_1__leaf_i_clk _0018_ VSS VSS VCC VCC instruction\[2\] sky130_fd_sc_hs__dfxtp_4
X_0912_ i_instruction[3] _0250_ _0273_ i_instruction[8] VSS VSS VCC VCC _0418_
+ sky130_fd_sc_hs__a22o_1
X_0843_ i_instruction[19] _0229_ _0195_ _0168_ VSS VSS VCC VCC _0357_ sky130_fd_sc_hs__a31o_1
X_0774_ _0177_ _0228_ _0260_ _0283_ VSS VSS VCC VCC _0296_ sky130_fd_sc_hs__or4_1
Xclkbuf_2_0_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_0_0_i_clk sky130_fd_sc_hs__clkbuf_8
X_0490_ o_csr_imm[0] _0086_ VSS VSS VCC VCC _0087_ sky130_fd_sc_hs__and2_1
X_1042_ o_csr_pc_next[5] VSS VSS VCC VCC o_pc_next[5] sky130_fd_sc_hs__buf_2
X_0826_ i_instruction[9] _0322_ VSS VSS VCC VCC _0342_ sky130_fd_sc_hs__and2_1
X_0757_ i_instruction[9] _0194_ _0273_ i_instruction[6] VSS VSS VCC VCC _0281_
+ sky130_fd_sc_hs__a22o_1
X_0688_ _0166_ instruction\[2\] _0167_ _0218_ VSS VSS VCC VCC _0018_ sky130_fd_sc_hs__o211a_1
X_0611_ o_csr_pc_next[7] i_pc_next[7] _0147_ VSS VSS VCC VCC _0154_ sky130_fd_sc_hs__mux2_1
X_0542_ o_funct3[0] _0095_ _0120_ VSS VSS VCC VCC o_imm_i[12] sky130_fd_sc_hs__a21o_2
X_0473_ instruction\[4\] _0074_ VSS VSS VCC VCC _0075_ sky130_fd_sc_hs__nor2_2
X_1025_ clknet_3_5__leaf_i_clk _0054_ VSS VSS VCC VCC o_pc[7] sky130_fd_sc_hs__dfxtp_2
X_0809_ _0249_ _0221_ _0315_ VSS VSS VCC VCC _0327_ sky130_fd_sc_hs__o21a_1
X_0525_ _0110_ VSS VSS VCC VCC o_imm_i[5] sky130_fd_sc_hs__buf_2
X_1008_ clknet_3_4__leaf_i_clk _0037_ VSS VSS VCC VCC o_csr_idx[1] sky130_fd_sc_hs__dfxtp_4
X_0508_ _0098_ VSS VSS VCC VCC _0099_ sky130_fd_sc_hs__buf_8
X_0790_ _0234_ _0200_ VSS VSS VCC VCC _0310_ sky130_fd_sc_hs__nor2_1
X_0988_ clknet_3_1__leaf_i_clk _0017_ VSS VSS VCC VCC instruction\[1\] sky130_fd_sc_hs__dfxtp_1
X_0911_ _0401_ _0416_ _0402_ VSS VSS VCC VCC _0417_ sky130_fd_sc_hs__o21a_1
X_0842_ _0353_ _0355_ _0289_ VSS VSS VCC VCC _0356_ sky130_fd_sc_hs__o21a_1
X_0773_ _0171_ i_instruction[11] VSS VSS VCC VCC _0295_ sky130_fd_sc_hs__and2_1
X_1041_ o_csr_pc_next[4] VSS VSS VCC VCC o_pc_next[4] sky130_fd_sc_hs__buf_2
X_0825_ _0211_ _0183_ _0184_ _0212_ VSS VSS VCC VCC _0341_ sky130_fd_sc_hs__o211a_4
X_0756_ _0251_ _0274_ _0198_ VSS VSS VCC VCC _0280_ sky130_fd_sc_hs__a21oi_1
X_0687_ _0195_ _0197_ _0205_ _0217_ VSS VSS VCC VCC _0218_ sky130_fd_sc_hs__a31o_1
X_0610_ _0153_ VSS VSS VCC VCC _0005_ sky130_fd_sc_hs__clkbuf_1
X_0541_ _0119_ VSS VSS VCC VCC _0120_ sky130_fd_sc_hs__buf_8
X_0472_ instruction\[6\] instruction\[3\] VSS VSS VCC VCC _0074_ sky130_fd_sc_hs__or2_2
X_1024_ clknet_3_0__leaf_i_clk _0053_ VSS VSS VCC VCC o_pc[6] sky130_fd_sc_hs__dfxtp_2
X_0808_ _0249_ _0325_ _0305_ VSS VSS VCC VCC _0326_ sky130_fd_sc_hs__a21o_1
X_0739_ _0229_ _0253_ _0264_ _0241_ VSS VSS VCC VCC _0265_ sky130_fd_sc_hs__a211o_1
X_0524_ o_csr_idx[5] _0085_ VSS VSS VCC VCC _0110_ sky130_fd_sc_hs__and2_1
X_1007_ clknet_3_4__leaf_i_clk _0036_ VSS VSS VCC VCC o_csr_idx[0] sky130_fd_sc_hs__dfxtp_4
X_0507_ _0096_ _0097_ VSS VSS VCC VCC _0098_ sky130_fd_sc_hs__and2_1
X_0987_ clknet_3_1__leaf_i_clk _0016_ VSS VSS VCC VCC instruction\[0\] sky130_fd_sc_hs__dfxtp_1
X_0910_ _0375_ _0224_ _0333_ i_instruction[3] VSS VSS VCC VCC _0416_ sky130_fd_sc_hs__a2bb2o_1
X_0841_ i_instruction[19] _0233_ _0331_ _0354_ VSS VSS VCC VCC _0355_ sky130_fd_sc_hs__a22o_1
X_0772_ _0166_ o_rd[3] _0167_ _0294_ VSS VSS VCC VCC _0026_ sky130_fd_sc_hs__o211a_1
X_1040_ o_csr_pc_next[3] VSS VSS VCC VCC o_pc_next[3] sky130_fd_sc_hs__buf_2
X_0824_ _0305_ _0284_ _0325_ i_instruction[9] VSS VSS VCC VCC _0340_ sky130_fd_sc_hs__a22o_1
X_0755_ _0243_ o_rd[1] _0267_ _0279_ _0248_ VSS VSS VCC VCC _0024_ sky130_fd_sc_hs__o221a_1
X_0686_ i_instruction[2] _0208_ _0210_ _0213_ _0216_ VSS VSS VCC VCC _0217_
+ sky130_fd_sc_hs__a221o_1
X_0540_ _0092_ _0118_ VSS VSS VCC VCC _0119_ sky130_fd_sc_hs__and2b_1
X_0471_ _0073_ VSS VSS VCC VCC o_op2_src sky130_fd_sc_hs__buf_2
X_1023_ clknet_3_5__leaf_i_clk _0052_ VSS VSS VCC VCC o_pc[5] sky130_fd_sc_hs__dfxtp_2
X_0807_ _0203_ _0201_ _0275_ VSS VSS VCC VCC _0325_ sky130_fd_sc_hs__a21oi_2
X_0738_ _0197_ _0258_ _0259_ _0263_ VSS VSS VCC VCC _0264_ sky130_fd_sc_hs__a31o_1
X_0669_ _0170_ i_instruction[3] VSS VSS VCC VCC _0200_ sky130_fd_sc_hs__nand2_4
X_0523_ _0108_ _0099_ _0109_ VSS VSS VCC VCC o_imm_i[4] sky130_fd_sc_hs__a21oi_4
X_1006_ clknet_3_6__leaf_i_clk _0035_ VSS VSS VCC VCC o_csr_imm[4] sky130_fd_sc_hs__dfxtp_4
X_0506_ o_inst_branch _0076_ VSS VSS VCC VCC _0097_ sky130_fd_sc_hs__nand2_1
X_0986_ clknet_3_1__leaf_i_clk _0015_ VSS VSS VCC VCC valid_input sky130_fd_sc_hs__dfxtp_1
X_0840_ i_instruction[11] _0221_ _0196_ VSS VSS VCC VCC _0354_ sky130_fd_sc_hs__and3_1
X_0771_ _0290_ _0293_ _0174_ VSS VSS VCC VCC _0294_ sky130_fd_sc_hs__a21o_1
X_0969_ o_pc[15] i_pc[15] _0446_ VSS VSS VCC VCC _0456_ sky130_fd_sc_hs__mux2_1
Xclkbuf_3_6__f_i_clk clknet_2_3_0_i_clk VSS VSS VCC VCC clknet_3_6__leaf_i_clk
+ sky130_fd_sc_hs__clkbuf_16
X_0823_ _0166_ o_csr_imm[1] _0309_ _0339_ VSS VSS VCC VCC _0032_ sky130_fd_sc_hs__o211a_1
X_0754_ _0229_ _0269_ _0272_ _0278_ VSS VSS VCC VCC _0279_ sky130_fd_sc_hs__a22o_1
X_0685_ _0210_ _0215_ i_stall VSS VSS VCC VCC _0216_ sky130_fd_sc_hs__a21o_1
X_0470_ o_inst_branch _0070_ _0072_ VSS VSS VCC VCC _0073_ sky130_fd_sc_hs__and3b_1
X_1022_ clknet_3_2__leaf_i_clk _0051_ VSS VSS VCC VCC o_pc[4] sky130_fd_sc_hs__dfxtp_2
X_0806_ _0321_ _0323_ _0261_ VSS VSS VCC VCC _0324_ sky130_fd_sc_hs__o21a_1
X_0737_ _0249_ _0232_ _0261_ _0262_ VSS VSS VCC VCC _0263_ sky130_fd_sc_hs__a22o_1
X_0668_ _0170_ i_instruction[2] VSS VSS VCC VCC _0199_ sky130_fd_sc_hs__nand2_4
X_0599_ o_csr_pc_next[1] i_pc_next[1] _0147_ VSS VSS VCC VCC _0148_ sky130_fd_sc_hs__mux2_1
X_0522_ o_rd[4] _0099_ _0086_ VSS VSS VCC VCC _0109_ sky130_fd_sc_hs__o21ai_1
X_1005_ clknet_3_1__leaf_i_clk _0034_ VSS VSS VCC VCC o_csr_imm[3] sky130_fd_sc_hs__dfxtp_2
X_0505_ _0096_ VSS VSS VCC VCC o_inst_store sky130_fd_sc_hs__inv_2

