* NGSPICE file created from rv_alu2.ext - technology: sky130A


X_3155_ _0805_ _0795_ net614 VSS VSS VCC VCC _1113_ sky130_fd_sc_hd__mux2_1
X_3086_ net620 _0904_ VSS VSS VCC VCC _1048_ sky130_fd_sc_hd__nor2_1
X_3988_ net515 net728 u_adder.i_cmp_inverse VSS VSS VCC VCC _1718_ sky130_fd_sc_hd__a21boi_1
X_2939_ net609 net409 VSS VSS VCC VCC _0909_ sky130_fd_sc_hd__nor2_4
X_4609_ _1869_ _1846_ _1845_ VSS VSS VCC VCC _2169_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_120_i_clk clknet_4_11__leaf_i_clk VSS VSS VCC VCC clknet_leaf_120_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_135_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_135_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4960_ _0928_ net400 VSS VSS VCC VCC _0404_ sky130_fd_sc_hd__nor2_1
X_3911_ u_pc_sel.i_pc_next\[2\] net116 net393 VSS VSS VCC VCC _0077_ sky130_fd_sc_hd__mux2_1
X_4891_ net479 _2425_ _2426_ net323 VSS VSS VCC VCC _2427_ sky130_fd_sc_hd__a31o_1
X_3842_ u_bits.i_op2\[14\] net726 _1663_ _1662_ VSS VSS VCC VCC _0058_ sky130_fd_sc_hd__o22a_1
X_3773_ net504 net236 net724 _1614_ VSS VSS VCC VCC _0038_ sky130_fd_sc_hd__o211a_1
X_2724_ net518 net525 _0696_ _0697_ VSS VSS VCC VCC _0699_ sky130_fd_sc_hd__a2bb2o_1
X_2655_ _0629_ _0627_ VSS VSS VCC VCC _0630_ sky130_fd_sc_hd__nand2_2
X_5374_ clknet_leaf_70_i_clk _0401_ VSS VSS VCC VCC u_muldiv.mul\[53\] sky130_fd_sc_hd__dfxtp_2
X_2586_ _0555_ _0558_ VSS VSS VCC VCC _0561_ sky130_fd_sc_hd__nand2_1
X_4325_ _1951_ _1952_ VSS VSS VCC VCC _1953_ sky130_fd_sc_hd__nand2_1
X_4256_ _1874_ _1881_ _1883_ VSS VSS VCC VCC _1884_ sky130_fd_sc_hd__a21oi_4
X_3207_ _1158_ _1160_ op_cnt\[0\] net39 _0432_ VSS VSS VCC VCC _0000_ sky130_fd_sc_hd__a2111oi_1
X_4187_ u_muldiv.mul\[17\] u_muldiv.mul\[16\] net404 VSS VSS VCC VCC _0231_
+ sky130_fd_sc_hd__mux2_1
X_3138_ _1030_ _1069_ VSS VSS VCC VCC _1097_ sky130_fd_sc_hd__or2_1
X_3069_ _0877_ _0927_ _1031_ VSS VSS VCC VCC _1032_ sky130_fd_sc_hd__nand3_2
Xfanout650 net651 VSS VSS VCC VCC net650 sky130_fd_sc_hd__buf_4
Xfanout661 u_bits.i_op1\[26\] VSS VSS VCC VCC net661 sky130_fd_sc_hd__clkbuf_4
Xfanout672 net673 VSS VSS VCC VCC net672 sky130_fd_sc_hd__buf_4
Xfanout683 u_bits.i_op1\[17\] VSS VSS VCC VCC net683 sky130_fd_sc_hd__clkbuf_16
Xfanout694 u_bits.i_op1\[12\] VSS VSS VCC VCC net694 sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_52_i_clk clknet_4_7__leaf_i_clk VSS VSS VCC VCC clknet_leaf_52_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_67_i_clk clknet_4_12__leaf_i_clk VSS VSS VCC VCC clknet_leaf_67_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2440_ u_muldiv.divisor\[13\] VSS VSS VCC VCC _0415_ sky130_fd_sc_hd__inv_2
X_4110_ net584 _1813_ net384 VSS VSS VCC VCC _1814_ sky130_fd_sc_hd__o21ai_1
X_5090_ clknet_leaf_73_i_clk _0123_ VSS VSS VCC VCC net306 sky130_fd_sc_hd__dfxtp_4
X_4041_ u_muldiv.divisor\[41\] net484 net335 u_muldiv.divisor\[42\] _1759_ vssd1 vssd1
+ vccd1 vccd1 _0161_ sky130_fd_sc_hd__a221o_1
X_4943_ _1183_ net402 VSS VSS VCC VCC _0387_ sky130_fd_sc_hd__nor2_1
X_4874_ _1973_ _2410_ net459 net479 VSS VSS VCC VCC _2411_ sky130_fd_sc_hd__a211o_1
X_3825_ net501 net78 net720 VSS VSS VCC VCC _1651_ sky130_fd_sc_hd__a21o_1
X_3756_ net671 net59 net389 VSS VSS VCC VCC _0025_ sky130_fd_sc_hd__mux2_1
X_2707_ _0674_ _0676_ _0678_ VSS VSS VCC VCC _0682_ sky130_fd_sc_hd__nand3b_2
X_3687_ net192 net354 net530 _1566_ VSS VSS VCC VCC _1567_ sky130_fd_sc_hd__a211o_1
X_2638_ net705 u_muldiv.add_prev\[7\] net540 VSS VSS VCC VCC _0613_ sky130_fd_sc_hd__mux2_2
Xoutput220 net220 VSS VSS VCC VCC o_pc_target[10] sky130_fd_sc_hd__buf_2
Xoutput231 net231 VSS VSS VCC VCC o_pc_target[6] sky130_fd_sc_hd__buf_2
Xoutput242 net242 VSS VSS VCC VCC o_res_src[0] sky130_fd_sc_hd__buf_2
Xoutput253 net253 VSS VSS VCC VCC o_result[17] sky130_fd_sc_hd__buf_2
Xoutput264 net264 VSS VSS VCC VCC o_result[27] sky130_fd_sc_hd__buf_2
X_5357_ clknet_leaf_103_i_clk _0384_ VSS VSS VCC VCC u_muldiv.mul\[36\] sky130_fd_sc_hd__dfxtp_1
Xoutput275 net275 VSS VSS VCC VCC o_result[8] sky130_fd_sc_hd__buf_2
X_2569_ _0537_ _0540_ net428 VSS VSS VCC VCC _0544_ sky130_fd_sc_hd__a21oi_2
Xoutput286 net286 VSS VSS VCC VCC o_wdata[16] sky130_fd_sc_hd__buf_2
Xoutput297 net297 VSS VSS VCC VCC o_wdata[26] sky130_fd_sc_hd__buf_2
X_4308_ _1934_ _1935_ VSS VSS VCC VCC _1936_ sky130_fd_sc_hd__or2_1
X_5288_ clknet_4_14__leaf_i_clk _0316_ VSS VSS VCC VCC u_muldiv.dividend\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_4239_ u_muldiv.divisor\[6\] u_muldiv.dividend\[6\] VSS VSS VCC VCC _1867_
+ sky130_fd_sc_hd__xnor2_2
Xfanout480 net481 VSS VSS VCC VCC net480 sky130_fd_sc_hd__clkbuf_4
Xfanout491 net495 VSS VSS VCC VCC net491 sky130_fd_sc_hd__clkbuf_4
X_3610_ _0932_ _1293_ _1294_ _1297_ net450 net455 VSS VSS VCC VCC _1495_ sky130_fd_sc_hd__mux4_1
X_4590_ _2150_ _2151_ net438 VSS VSS VCC VCC _2152_ sky130_fd_sc_hd__a21oi_1
X_3541_ net352 _1425_ _1429_ _1430_ VSS VSS VCC VCC _1431_ sky130_fd_sc_hd__a31o_1
X_3472_ net611 _1363_ _1364_ net604 VSS VSS VCC VCC _1366_ sky130_fd_sc_hd__o211ai_2
X_5211_ clknet_leaf_18_i_clk _0243_ VSS VSS VCC VCC u_muldiv.mul\[28\] sky130_fd_sc_hd__dfxtp_1
X_5142_ clknet_4_4__leaf_i_clk _0174_ VSS VSS VCC VCC u_muldiv.divisor\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_5073_ clknet_leaf_78_i_clk _0106_ VSS VSS VCC VCC net223 sky130_fd_sc_hd__dfxtp_1
X_4024_ net600 net599 _1737_ net379 VSS VSS VCC VCC _1746_ sky130_fd_sc_hd__o31a_1
X_4926_ _1146_ _2428_ _2429_ VSS VSS VCC VCC _2430_ sky130_fd_sc_hd__and3_1
X_4857_ _2394_ _2395_ net476 VSS VSS VCC VCC _2396_ sky130_fd_sc_hd__o21a_1
X_3808_ net506 _1637_ VSS VSS VCC VCC _1638_ sky130_fd_sc_hd__and2b_1
X_4788_ _2322_ u_muldiv.dividend\[22\] net434 VSS VSS VCC VCC _2333_ sky130_fd_sc_hd__a21o_1
X_3739_ u_bits.i_op1\[5\] net72 net389 VSS VSS VCC VCC _0008_ sky130_fd_sc_hd__mux2_1
X_2972_ net454 _0937_ _0939_ VSS VSS VCC VCC _0940_ sky130_fd_sc_hd__o21ai_1
X_4711_ u_muldiv.dividend\[15\] u_muldiv.dividend\[14\] u_muldiv.dividend\[16\] _2239_
+ VSS VSS VCC VCC _2262_ sky130_fd_sc_hd__or4_4
X_4642_ u_muldiv.dividend\[9\] net324 net375 _2199_ VSS VSS VCC VCC _0322_
+ sky130_fd_sc_hd__a31o_1
X_4573_ u_muldiv.dividend\[0\] net464 u_muldiv.dividend\[3\] net463 vssd1 vssd1 vccd1
+ vccd1 _2137_ sky130_fd_sc_hd__or4_1
X_3524_ net617 _0910_ _0850_ net353 _1414_ VSS VSS VCC VCC _1415_ sky130_fd_sc_hd__o311a_1
X_3455_ _1346_ net367 net572 _1349_ VSS VSS VCC VCC _1350_ sky130_fd_sc_hd__a31o_1
X_3386_ net359 net183 _1282_ _1283_ VSS VSS VCC VCC _1284_ sky130_fd_sc_hd__a211o_1
X_5125_ clknet_leaf_28_i_clk _0157_ VSS VSS VCC VCC u_muldiv.divisor\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_5056_ clknet_leaf_34_i_clk _0089_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_4007_ _1732_ net383 _1731_ VSS VSS VCC VCC _1733_ sky130_fd_sc_hd__and3b_1
X_4909_ u_muldiv.divisor\[16\] net488 net341 u_muldiv.divisor\[17\] vssd1 vssd1 vccd1
+ vccd1 _0361_ sky130_fd_sc_hd__a22o_1
X_3240_ _0630_ _0605_ _0727_ _0635_ VSS VSS VCC VCC _1184_ sky130_fd_sc_hd__o211a_1
X_3171_ net651 u_muldiv.add_prev\[31\] net532 VSS VSS VCC VCC _1128_ sky130_fd_sc_hd__mux2_1
X_2955_ _0922_ _0923_ VSS VSS VCC VCC _0924_ sky130_fd_sc_hd__and2_1
X_2886_ net669 net674 net671 net675 net634 net639 VSS VSS VCC VCC _0858_ sky130_fd_sc_hd__mux4_1
X_4625_ _2143_ _2171_ _0435_ _0436_ VSS VSS VCC VCC _2184_ sky130_fd_sc_hd__nand4_2
X_4556_ _1855_ _1856_ _1858_ _1860_ _2120_ VSS VSS VCC VCC _2121_ sky130_fd_sc_hd__a41o_1
X_3507_ net607 net614 _0815_ _0795_ VSS VSS VCC VCC _1399_ sky130_fd_sc_hd__or4_1
X_4487_ net465 u_muldiv.quotient_msk\[26\] net433 _2088_ _2089_ vssd1 vssd1 vccd1
+ vccd1 _2090_ sky130_fd_sc_hd__a32o_1
X_3438_ net557 u_muldiv.mul\[2\] net414 net529 _1333_ VSS VSS VCC VCC _1334_
+ sky130_fd_sc_hd__o311a_1
X_3369_ _1242_ _1266_ VSS VSS VCC VCC _1267_ sky130_fd_sc_hd__nand2_1
X_5108_ clknet_leaf_8_i_clk _0141_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_5039_ clknet_leaf_44_i_clk _0072_ VSS VSS VCC VCC u_bits.i_op2\[28\] sky130_fd_sc_hd__dfxtp_4
Xinput120 i_pc_next[6] VSS VSS VCC VCC net120 sky130_fd_sc_hd__clkbuf_2
Xinput131 i_pc_target[2] VSS VSS VCC VCC net131 sky130_fd_sc_hd__buf_2
Xinput142 i_rd[3] VSS VSS VCC VCC net142 sky130_fd_sc_hd__clkbuf_2
Xinput153 i_reg_data2[18] VSS VSS VCC VCC net153 sky130_fd_sc_hd__clkbuf_1
Xinput164 i_reg_data2[28] VSS VSS VCC VCC net164 sky130_fd_sc_hd__clkbuf_1
Xinput175 i_reg_data2[9] VSS VSS VCC VCC net175 sky130_fd_sc_hd__clkbuf_1
X_2740_ _0713_ _0714_ VSS VSS VCC VCC _0715_ sky130_fd_sc_hd__nand2_1
X_2671_ _0642_ _0643_ _0645_ VSS VSS VCC VCC _0646_ sky130_fd_sc_hd__nand3_4
X_4410_ u_muldiv.o_div\[9\] _2020_ u_muldiv.o_div\[10\] VSS VSS VCC VCC _2029_
+ sky130_fd_sc_hd__o21ai_1
X_4341_ _1967_ _1960_ _1968_ VSS VSS VCC VCC _1969_ sky130_fd_sc_hd__o21ai_2
X_4272_ _0415_ u_muldiv.dividend\[13\] _1899_ VSS VSS VCC VCC _1900_ sky130_fd_sc_hd__a21bo_1
X_3223_ _0606_ _0629_ _0633_ VSS VSS VCC VCC _1171_ sky130_fd_sc_hd__a21oi_2
X_3154_ u_muldiv.mul\[62\] net363 net357 u_muldiv.mul\[30\] VSS VSS VCC VCC
+ _1112_ sky130_fd_sc_hd__a22o_1
X_3085_ net451 _1044_ _1046_ VSS VSS VCC VCC _1047_ sky130_fd_sc_hd__o21ai_4
X_3987_ u_wr_mux.i_reg_data2\[31\] net168 net396 VSS VSS VCC VCC _0149_ sky130_fd_sc_hd__mux2_1
X_2938_ net453 net450 VSS VSS VCC VCC _0908_ sky130_fd_sc_hd__nand2_4
X_2869_ u_bits.i_sra net458 net650 _0774_ VSS VSS VCC VCC _0841_ sky130_fd_sc_hd__o211a_1
X_4608_ u_muldiv.dividend\[6\] net325 net376 _2168_ VSS VSS VCC VCC _0319_
+ sky130_fd_sc_hd__a31o_1
X_4539_ u_muldiv.quotient_msk\[27\] net476 net332 u_muldiv.quotient_msk\[28\] vssd1
+ vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__a22o_1
X_3910_ u_pc_sel.i_pc_next\[1\] net115 net388 VSS VSS VCC VCC _0076_ sky130_fd_sc_hd__mux2_1
X_4890_ u_muldiv.dividend\[31\] _2412_ VSS VSS VCC VCC _2426_ sky130_fd_sc_hd__or2_1
X_3841_ net508 net82 net719 VSS VSS VCC VCC _1663_ sky130_fd_sc_hd__a21o_1
X_3772_ net140 net504 VSS VSS VCC VCC _1614_ sky130_fd_sc_hd__nand2b_1
X_2723_ _0697_ _0457_ _0696_ VSS VSS VCC VCC _0698_ sky130_fd_sc_hd__nand3_1
X_2654_ _0591_ _0599_ _0601_ VSS VSS VCC VCC _0629_ sky130_fd_sc_hd__o21a_1
X_5373_ clknet_leaf_151_i_clk _0400_ VSS VSS VCC VCC u_muldiv.mul\[52\] sky130_fd_sc_hd__dfxtp_1
X_2585_ _0556_ _0557_ _0552_ _0553_ VSS VSS VCC VCC _0560_ sky130_fd_sc_hd__o211ai_4
X_4324_ _0448_ u_muldiv.divisor\[27\] VSS VSS VCC VCC _1952_ sky130_fd_sc_hd__nand2_1
X_4255_ u_muldiv.divisor\[8\] _1882_ _1880_ VSS VSS VCC VCC _1883_ sky130_fd_sc_hd__o21ai_1
X_3206_ _1158_ _1160_ op_cnt\[0\] VSS VSS VCC VCC _1161_ sky130_fd_sc_hd__a21oi_2
X_4186_ u_muldiv.mul\[16\] u_muldiv.mul\[15\] net404 VSS VSS VCC VCC _0230_
+ sky130_fd_sc_hd__mux2_1
X_3137_ net731 net27 _1096_ VSS VSS VCC VCC net266 sky130_fd_sc_hd__o21a_1
X_3068_ _0964_ _0965_ _0997_ _0998_ VSS VSS VCC VCC _1031_ sky130_fd_sc_hd__and4_1
Xfanout640 net641 VSS VSS VCC VCC net640 sky130_fd_sc_hd__buf_4
Xfanout651 u_bits.i_op1\[31\] VSS VSS VCC VCC net651 sky130_fd_sc_hd__clkbuf_8
Xfanout662 net663 VSS VSS VCC VCC net662 sky130_fd_sc_hd__buf_4
Xfanout673 net674 VSS VSS VCC VCC net673 sky130_fd_sc_hd__buf_4
Xfanout684 net685 VSS VSS VCC VCC net684 sky130_fd_sc_hd__clkbuf_4
Xfanout695 u_bits.i_op1\[11\] VSS VSS VCC VCC net695 sky130_fd_sc_hd__buf_6
X_4040_ net595 _1757_ _1758_ VSS VSS VCC VCC _1759_ sky130_fd_sc_hd__o21ba_1
X_4942_ _1173_ _1174_ net407 VSS VSS VCC VCC _0386_ sky130_fd_sc_hd__and3_1
X_4873_ _1967_ _1960_ _2409_ VSS VSS VCC VCC _2410_ sky130_fd_sc_hd__o21ai_1
X_3824_ net503 _1649_ VSS VSS VCC VCC _1650_ sky130_fd_sc_hd__and2b_1
X_3755_ net673 net58 net394 VSS VSS VCC VCC _0024_ sky130_fd_sc_hd__mux2_1
X_2706_ _0674_ _0677_ _0675_ VSS VSS VCC VCC _0681_ sky130_fd_sc_hd__nor3_2
X_3686_ _1561_ _1565_ net522 VSS VSS VCC VCC _1566_ sky130_fd_sc_hd__o21ba_1
Xoutput210 net210 VSS VSS VCC VCC o_add[5] sky130_fd_sc_hd__buf_2
X_2637_ _0608_ _0457_ VSS VSS VCC VCC _0612_ sky130_fd_sc_hd__nand2_1
Xoutput221 net221 VSS VSS VCC VCC o_pc_target[11] sky130_fd_sc_hd__buf_2
Xoutput232 net232 VSS VSS VCC VCC o_pc_target[7] sky130_fd_sc_hd__buf_2
Xoutput243 net577 VSS VSS VCC VCC o_res_src[1] sky130_fd_sc_hd__buf_2
Xoutput254 net254 VSS VSS VCC VCC o_result[18] sky130_fd_sc_hd__buf_2
X_5356_ clknet_leaf_100_i_clk _0383_ VSS VSS VCC VCC u_muldiv.mul\[35\] sky130_fd_sc_hd__dfxtp_1
X_2568_ net518 net525 _0541_ VSS VSS VCC VCC _0543_ sky130_fd_sc_hd__o21ai_1
Xoutput265 net265 VSS VSS VCC VCC o_result[28] sky130_fd_sc_hd__buf_2
Xoutput276 net276 VSS VSS VCC VCC o_result[9] sky130_fd_sc_hd__buf_2
Xoutput287 net287 VSS VSS VCC VCC o_wdata[17] sky130_fd_sc_hd__buf_2
Xoutput298 net298 VSS VSS VCC VCC o_wdata[27] sky130_fd_sc_hd__buf_2
X_4307_ u_muldiv.dividend\[20\] u_muldiv.divisor\[20\] VSS VSS VCC VCC _1935_
+ sky130_fd_sc_hd__and2b_1
X_5287_ clknet_leaf_87_i_clk _0315_ VSS VSS VCC VCC u_muldiv.dividend\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2499_ _0470_ _0472_ VSS VSS VCC VCC _0474_ sky130_fd_sc_hd__nand2_1
X_4238_ _1865_ _1849_ _1850_ _1847_ VSS VSS VCC VCC _1866_ sky130_fd_sc_hd__a31oi_4
X_4169_ net550 net499 net206 VSS VSS VCC VCC _0213_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_134_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_134_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout470 net472 VSS VSS VCC VCC net470 sky130_fd_sc_hd__buf_6
Xfanout481 net487 VSS VSS VCC VCC net481 sky130_fd_sc_hd__buf_4
Xfanout492 net494 VSS VSS VCC VCC net492 sky130_fd_sc_hd__buf_4
X_3540_ u_bits.i_op2\[8\] net702 net352 VSS VSS VCC VCC _1430_ sky130_fd_sc_hd__a21oi_1
X_3471_ net612 _1363_ _1364_ VSS VSS VCC VCC _1365_ sky130_fd_sc_hd__o21ai_1
X_5210_ clknet_leaf_156_i_clk _0242_ VSS VSS VCC VCC u_muldiv.mul\[27\] sky130_fd_sc_hd__dfxtp_1
X_5141_ clknet_leaf_36_i_clk _0173_ VSS VSS VCC VCC u_muldiv.divisor\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_5072_ clknet_leaf_135_i_clk _0105_ VSS VSS VCC VCC net222 sky130_fd_sc_hd__dfxtp_1
X_4023_ net603 net600 net599 _1279_ VSS VSS VCC VCC _1745_ sky130_fd_sc_hd__or4_1
X_4925_ u_bits.i_op1\[31\] net579 net416 VSS VSS VCC VCC _2429_ sky130_fd_sc_hd__o21a_1
X_4856_ u_muldiv.dividend\[27\] u_muldiv.dividend\[26\] u_muldiv.dividend\[25\] _2345_
+ u_muldiv.dividend\[28\] VSS VSS VCC VCC _2395_ sky130_fd_sc_hd__o41a_1
X_3807_ net598 net600 net546 VSS VSS VCC VCC _1637_ sky130_fd_sc_hd__mux2_1
X_4787_ net467 _2330_ _2331_ _2328_ VSS VSS VCC VCC _2332_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_51_i_clk clknet_4_7__leaf_i_clk VSS VSS VCC VCC clknet_leaf_51_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3738_ net711 net71 net398 VSS VSS VCC VCC _0007_ sky130_fd_sc_hd__mux2_1
X_3669_ _0429_ net569 net683 VSS VSS VCC VCC _1550_ sky130_fd_sc_hd__or3b_1
X_5339_ clknet_leaf_166_i_clk _0367_ VSS VSS VCC VCC u_muldiv.divisor\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_19_i_clk clknet_4_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_19_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2971_ net620 _0938_ VSS VSS VCC VCC _0939_ sky130_fd_sc_hd__or2_1
X_4710_ _2258_ u_muldiv.dividend\[16\] VSS VSS VCC VCC _2261_ sky130_fd_sc_hd__nand2_1
X_4641_ _2192_ _2198_ net322 VSS VSS VCC VCC _2199_ sky130_fd_sc_hd__a21oi_1
X_4572_ u_muldiv.dividend\[0\] net464 u_muldiv.dividend\[3\] net463 vssd1 vssd1 vccd1
+ vccd1 _2136_ sky130_fd_sc_hd__nor4_4
X_3523_ u_bits.i_op2\[7\] net705 net351 _1413_ VSS VSS VCC VCC _1414_ sky130_fd_sc_hd__o211ai_1
X_3454_ _0848_ _0907_ _0909_ _1348_ net412 VSS VSS VCC VCC _1349_ sky130_fd_sc_hd__a311o_1
X_3385_ _0896_ _0907_ net345 net412 VSS VSS VCC VCC _1283_ sky130_fd_sc_hd__a31o_1
X_5124_ clknet_leaf_28_i_clk _0156_ VSS VSS VCC VCC u_muldiv.divisor\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_5055_ clknet_leaf_61_i_clk _0088_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[13\]
+ sky130_fd_sc_hd__dfxtp_4
X_4006_ net640 net626 net624 net618 net378 VSS VSS VCC VCC _1732_ sky130_fd_sc_hd__o311a_1
X_4908_ u_muldiv.divisor\[15\] net489 net341 u_muldiv.divisor\[16\] vssd1 vssd1 vccd1
+ vccd1 _0360_ sky130_fd_sc_hd__a22o_1
X_4839_ net667 net664 net662 net660 VSS VSS VCC VCC _2379_ sky130_fd_sc_hd__nor4_1
X_3170_ net577 _1127_ VSS VSS VCC VCC net268 sky130_fd_sc_hd__and2b_1
X_2954_ net663 u_muldiv.add_prev\[25\] net534 VSS VSS VCC VCC _0923_ sky130_fd_sc_hd__mux2_1
X_2885_ net604 net450 VSS VSS VCC VCC _0857_ sky130_fd_sc_hd__or2_1
X_4624_ _1876_ _1877_ _1874_ VSS VSS VCC VCC _2183_ sky130_fd_sc_hd__a21o_1
X_4555_ _2119_ net473 VSS VSS VCC VCC _2120_ sky130_fd_sc_hd__nand2_1
X_3506_ net606 _0779_ _0856_ _1395_ _1397_ VSS VSS VCC VCC _1398_ sky130_fd_sc_hd__a221o_1
X_4486_ u_muldiv.o_div\[25\] _2081_ u_muldiv.o_div\[26\] VSS VSS VCC VCC _2089_
+ sky130_fd_sc_hd__o21ai_1
X_3437_ u_muldiv.o_div\[2\] net366 net359 _1332_ VSS VSS VCC VCC _1333_ sky130_fd_sc_hd__a211o_1
X_3368_ net571 net560 VSS VSS VCC VCC _1266_ sky130_fd_sc_hd__and2b_1
X_5107_ clknet_leaf_48_i_clk _0140_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_3299_ _0753_ _1221_ _0889_ VSS VSS VCC VCC _1229_ sky130_fd_sc_hd__nand3_1
X_5038_ clknet_leaf_14_i_clk _0071_ VSS VSS VCC VCC u_bits.i_op2\[27\] sky130_fd_sc_hd__dfxtp_4
Xinput110 i_pc_next[11] VSS VSS VCC VCC net110 sky130_fd_sc_hd__clkbuf_1
Xinput121 i_pc_next[7] VSS VSS VCC VCC net121 sky130_fd_sc_hd__clkbuf_1
Xinput132 i_pc_target[3] VSS VSS VCC VCC net132 sky130_fd_sc_hd__buf_4
Xinput143 i_rd[4] VSS VSS VCC VCC net143 sky130_fd_sc_hd__clkbuf_1
Xinput154 i_reg_data2[19] VSS VSS VCC VCC net154 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput165 i_reg_data2[29] VSS VSS VCC VCC net165 sky130_fd_sc_hd__clkbuf_2
Xinput176 i_reg_write VSS VSS VCC VCC net176 sky130_fd_sc_hd__buf_6
X_2670_ net694 u_muldiv.add_prev\[12\] net542 VSS VSS VCC VCC _0645_ sky130_fd_sc_hd__mux2_1
X_4340_ _1963_ _1964_ _1961_ VSS VSS VCC VCC _1968_ sky130_fd_sc_hd__a21oi_1
X_4271_ _0415_ u_muldiv.dividend\[13\] _1895_ VSS VSS VCC VCC _1899_ sky130_fd_sc_hd__o21ai_1
X_3222_ _1170_ VSS VSS VCC VCC net209 sky130_fd_sc_hd__inv_6
X_3153_ u_muldiv.dividend\[30\] net419 net364 u_muldiv.o_div\[30\] net442 vssd1 vssd1
+ vccd1 vccd1 _1111_ sky130_fd_sc_hd__a221o_1
X_3084_ net613 _1045_ VSS VSS VCC VCC _1046_ sky130_fd_sc_hd__or2_1
X_3986_ u_wr_mux.i_reg_data2\[30\] net167 net387 VSS VSS VCC VCC _0148_ sky130_fd_sc_hd__mux2_1
X_2937_ net621 net614 VSS VSS VCC VCC _0907_ sky130_fd_sc_hd__nor2_4
X_2868_ net644 net634 VSS VSS VCC VCC _0840_ sky130_fd_sc_hd__nor2_2
X_4607_ net497 _2167_ _2162_ net320 VSS VSS VCC VCC _2168_ sky130_fd_sc_hd__o211a_1
X_2799_ net650 u_bits.i_sra net455 VSS VSS VCC VCC _0773_ sky130_fd_sc_hd__a21o_1
X_4538_ u_muldiv.quotient_msk\[26\] net475 net332 u_muldiv.quotient_msk\[27\] vssd1
+ vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__a22o_1
X_4469_ u_muldiv.quotient_msk\[22\] u_muldiv.o_div\[22\] net469 net437 vssd1 vssd1
+ vccd1 vccd1 _2076_ sky130_fd_sc_hd__o211a_1
X_3840_ net508 _1661_ VSS VSS VCC VCC _1662_ sky130_fd_sc_hd__and2b_1
X_3771_ net514 net235 net727 _1613_ VSS VSS VCC VCC _0037_ sky130_fd_sc_hd__o211a_1
X_2722_ net648 net554 net696 net542 net425 VSS VSS VCC VCC _0697_ sky130_fd_sc_hd__o2111ai_4
X_2653_ _0591_ _0599_ _0601_ VSS VSS VCC VCC _0628_ sky130_fd_sc_hd__o21ai_2
X_2584_ _0556_ _0557_ _0552_ _0553_ VSS VSS VCC VCC _0559_ sky130_fd_sc_hd__o211a_1
X_5372_ clknet_leaf_151_i_clk _0399_ VSS VSS VCC VCC u_muldiv.mul\[51\] sky130_fd_sc_hd__dfxtp_1
X_4323_ u_muldiv.divisor\[27\] _0448_ VSS VSS VCC VCC _1951_ sky130_fd_sc_hd__or2_1
X_4254_ _1844_ u_muldiv.dividend\[8\] VSS VSS VCC VCC _1882_ sky130_fd_sc_hd__nand2_1
X_3205_ net548 op_cnt\[5\] _1159_ op_cnt\[4\] VSS VSS VCC VCC _1160_ sky130_fd_sc_hd__or4bb_1
X_4185_ u_muldiv.mul\[15\] u_muldiv.mul\[14\] net404 VSS VSS VCC VCC _0229_
+ sky130_fd_sc_hd__mux2_1
X_3136_ net577 _1095_ VSS VSS VCC VCC _1096_ sky130_fd_sc_hd__nor2_1
X_3067_ _1028_ _1029_ VSS VSS VCC VCC _1030_ sky130_fd_sc_hd__nand2_4
X_3969_ u_wr_mux.i_reg_data2\[13\] net148 net386 VSS VSS VCC VCC _0131_ sky130_fd_sc_hd__mux2_1
Xfanout630 net631 VSS VSS VCC VCC net630 sky130_fd_sc_hd__buf_4
Xfanout641 u_bits.i_op2\[0\] VSS VSS VCC VCC net641 sky130_fd_sc_hd__buf_8
Xfanout652 net653 VSS VSS VCC VCC net652 sky130_fd_sc_hd__buf_6
Xfanout663 u_bits.i_op1\[25\] VSS VSS VCC VCC net663 sky130_fd_sc_hd__buf_6
Xfanout674 u_bits.i_op1\[21\] VSS VSS VCC VCC net674 sky130_fd_sc_hd__buf_8
Xfanout685 u_bits.i_op1\[16\] VSS VSS VCC VCC net685 sky130_fd_sc_hd__buf_12
Xfanout696 u_bits.i_op1\[11\] VSS VSS VCC VCC net696 sky130_fd_sc_hd__buf_4
X_4941_ _1172_ _1176_ net406 VSS VSS VCC VCC _0385_ sky130_fd_sc_hd__and3_1
X_4872_ _1963_ _1964_ _1970_ _1971_ _1961_ VSS VSS VCC VCC _2409_ sky130_fd_sc_hd__a2111oi_1
X_3823_ net594 net596 net546 VSS VSS VCC VCC _1649_ sky130_fd_sc_hd__mux2_1
X_3754_ net675 net57 net393 VSS VSS VCC VCC _0023_ sky130_fd_sc_hd__mux2_1
X_2705_ _0674_ _0675_ _0677_ VSS VSS VCC VCC _0680_ sky130_fd_sc_hd__o21ai_2
X_3685_ net588 net680 net410 _1559_ _1564_ VSS VSS VCC VCC _1565_ sky130_fd_sc_hd__a311o_1
Xoutput200 net200 VSS VSS VCC VCC o_add[25] sky130_fd_sc_hd__buf_2
X_2636_ net540 _0426_ net518 net525 _0607_ VSS VSS VCC VCC _0611_ sky130_fd_sc_hd__o221ai_4
Xoutput211 net211 VSS VSS VCC VCC o_add[6] sky130_fd_sc_hd__buf_2
Xoutput222 net222 VSS VSS VCC VCC o_pc_target[12] sky130_fd_sc_hd__buf_2
Xoutput233 net233 VSS VSS VCC VCC o_pc_target[8] sky130_fd_sc_hd__buf_2
Xoutput244 net244 VSS VSS VCC VCC o_res_src[2] sky130_fd_sc_hd__buf_2
X_5355_ clknet_leaf_100_i_clk _0382_ VSS VSS VCC VCC u_muldiv.mul\[34\] sky130_fd_sc_hd__dfxtp_1
Xoutput255 net255 VSS VSS VCC VCC o_result[19] sky130_fd_sc_hd__buf_2
X_2567_ _0460_ _0539_ _0537_ net432 VSS VSS VCC VCC _0542_ sky130_fd_sc_hd__o211ai_2
Xoutput266 net266 VSS VSS VCC VCC o_result[29] sky130_fd_sc_hd__buf_2
Xoutput277 net277 VSS VSS VCC VCC o_store sky130_fd_sc_hd__buf_2
Xoutput288 net288 VSS VSS VCC VCC o_wdata[18] sky130_fd_sc_hd__buf_2
X_4306_ u_muldiv.divisor\[20\] u_muldiv.dividend\[20\] VSS VSS VCC VCC _1934_
+ sky130_fd_sc_hd__and2b_1
Xoutput299 net299 VSS VSS VCC VCC o_wdata[28] sky130_fd_sc_hd__buf_2
X_5286_ clknet_leaf_87_i_clk _0314_ VSS VSS VCC VCC u_muldiv.dividend\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2498_ _0470_ _0472_ VSS VSS VCC VCC _0473_ sky130_fd_sc_hd__and2_1
X_4237_ u_muldiv.divisor\[3\] _0441_ _1851_ _1863_ VSS VSS VCC VCC _1865_
+ sky130_fd_sc_hd__o211ai_4
X_4168_ _1071_ _1072_ net400 VSS VSS VCC VCC _0212_ sky130_fd_sc_hd__and3_1
X_3119_ net602 _1078_ net327 VSS VSS VCC VCC _1079_ sky130_fd_sc_hd__o21a_1
X_4099_ u_muldiv.divisor\[53\] net484 net335 u_muldiv.divisor\[54\] _1805_ vssd1 vssd1
+ vccd1 vccd1 _0173_ sky130_fd_sc_hd__a221o_1
Xfanout460 u_bits.i_op1\[0\] VSS VSS VCC VCC net460 sky130_fd_sc_hd__buf_4
Xfanout471 net472 VSS VSS VCC VCC net471 sky130_fd_sc_hd__buf_2
Xfanout482 net483 VSS VSS VCC VCC net482 sky130_fd_sc_hd__clkbuf_4
Xfanout493 net494 VSS VSS VCC VCC net493 sky130_fd_sc_hd__clkbuf_4
X_3470_ net612 _1039_ VSS VSS VCC VCC _1364_ sky130_fd_sc_hd__nand2_1
X_5140_ clknet_leaf_36_i_clk _0172_ VSS VSS VCC VCC u_muldiv.divisor\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_5071_ clknet_4_15__leaf_i_clk _0104_ VSS VSS VCC VCC net221 sky130_fd_sc_hd__dfxtp_4
X_4022_ u_muldiv.divisor\[37\] net482 net337 u_muldiv.divisor\[38\] _1744_ vssd1 vssd1
+ vccd1 vccd1 _0157_ sky130_fd_sc_hd__a221o_1
X_4924_ net581 net580 net579 _1827_ VSS VSS VCC VCC _2428_ sky130_fd_sc_hd__or4_1
X_4855_ u_muldiv.dividend\[28\] _2384_ VSS VSS VCC VCC _2394_ sky130_fd_sc_hd__nor2_1
X_3806_ net600 net724 _1636_ _1635_ VSS VSS VCC VCC _0049_ sky130_fd_sc_hd__o22a_1
X_4786_ net672 _2316_ net371 net670 VSS VSS VCC VCC _2331_ sky130_fd_sc_hd__o211a_1
X_3737_ net714 net70 net397 VSS VSS VCC VCC _0006_ sky130_fd_sc_hd__mux2_1
X_3668_ _0945_ _0806_ _0856_ _0940_ _1548_ VSS VSS VCC VCC _1549_ sky130_fd_sc_hd__a221o_1
X_2619_ net649 net554 net708 net539 net425 VSS VSS VCC VCC _0594_ sky130_fd_sc_hd__o2111ai_4
X_3599_ net573 net422 _1481_ net520 VSS VSS VCC VCC _1485_ sky130_fd_sc_hd__a31o_1
X_5338_ clknet_leaf_164_i_clk _0366_ VSS VSS VCC VCC u_muldiv.divisor\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_5269_ clknet_leaf_128_i_clk _0297_ VSS VSS VCC VCC u_muldiv.quotient_msk\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_2970_ net699 net701 net704 net706 net642 net630 VSS VSS VCC VCC _0938_ sky130_fd_sc_hd__mux4_1
X_4640_ net435 _2193_ _2194_ _2196_ _2197_ VSS VSS VCC VCC _2198_ sky130_fd_sc_hd__o32a_1
X_4571_ _2130_ net473 _2129_ _2134_ VSS VSS VCC VCC _2135_ sky130_fd_sc_hd__a31o_1
X_3522_ net566 _0436_ _0426_ VSS VSS VCC VCC _1413_ sky130_fd_sc_hd__or3_1
Xclkbuf_4_14__f_i_clk clknet_2_3_0_i_clk VSS VSS VCC VCC clknet_4_14__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3453_ net617 net712 net351 _1347_ VSS VSS VCC VCC _1348_ sky130_fd_sc_hd__o211a_1
X_3384_ net643 net460 _1281_ VSS VSS VCC VCC _1282_ sky130_fd_sc_hd__o21a_1
X_5123_ clknet_leaf_16_i_clk _0155_ VSS VSS VCC VCC u_muldiv.divisor\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_5054_ clknet_4_15__leaf_i_clk _0087_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[12\]
+ sky130_fd_sc_hd__dfxtp_4
X_4005_ net624 net378 _1728_ net618 VSS VSS VCC VCC _1731_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_133_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_133_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4907_ u_muldiv.divisor\[14\] net489 net341 u_muldiv.divisor\[15\] vssd1 vssd1 vccd1
+ vccd1 _0359_ sky130_fd_sc_hd__a22o_1
X_4838_ _1953_ _2376_ _2377_ VSS VSS VCC VCC _2378_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_148_i_clk clknet_4_8__leaf_i_clk VSS VSS VCC VCC clknet_leaf_148_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4769_ _1937_ _1939_ _2313_ VSS VSS VCC VCC _2315_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_50_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_50_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2953_ net427 _0921_ VSS VSS VCC VCC _0922_ sky130_fd_sc_hd__xor2_1
X_2884_ net608 net452 VSS VSS VCC VCC _0856_ sky130_fd_sc_hd__nor2_4
X_4623_ _2180_ _2181_ net435 VSS VSS VCC VCC _2182_ sky130_fd_sc_hd__a21o_1
X_4554_ _1855_ _1856_ _1858_ _1860_ VSS VSS VCC VCC _2119_ sky130_fd_sc_hd__a22o_1
X_3505_ net606 _1396_ _0765_ VSS VSS VCC VCC _1397_ sky130_fd_sc_hd__o21ai_1
X_4485_ u_muldiv.o_div\[25\] u_muldiv.o_div\[26\] _2081_ net475 vssd1 vssd1 vccd1
+ vccd1 _2088_ sky130_fd_sc_hd__o31a_1
X_3436_ net568 net557 net463 u_muldiv.mul\[34\] net361 VSS VSS VCC VCC _1332_
+ sky130_fd_sc_hd__a32o_1
X_3367_ net415 net183 net566 net194 VSS VSS VCC VCC net314 sky130_fd_sc_hd__o22a_2
X_5106_ clknet_leaf_119_i_clk _0139_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[21\]
+ sky130_fd_sc_hd__dfxtp_2
X_3298_ _1227_ _1188_ _1204_ _1196_ VSS VSS VCC VCC _1228_ sky130_fd_sc_hd__nand4_2
X_5037_ clknet_leaf_12_i_clk _0070_ VSS VSS VCC VCC u_bits.i_op2\[26\] sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_18_i_clk clknet_4_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_18_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput100 i_op2[30] VSS VSS VCC VCC net100 sky130_fd_sc_hd__clkbuf_8
Xinput111 i_pc_next[12] VSS VSS VCC VCC net111 sky130_fd_sc_hd__clkbuf_1
Xinput122 i_pc_next[8] VSS VSS VCC VCC net122 sky130_fd_sc_hd__clkbuf_4
Xinput133 i_pc_target[4] VSS VSS VCC VCC net133 sky130_fd_sc_hd__clkbuf_4
Xinput144 i_reg_data2[0] VSS VSS VCC VCC net144 sky130_fd_sc_hd__clkbuf_1
Xinput155 i_reg_data2[1] VSS VSS VCC VCC net155 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput166 i_reg_data2[2] VSS VSS VCC VCC net166 sky130_fd_sc_hd__clkbuf_1
Xinput177 i_res_src[0] VSS VSS VCC VCC net177 sky130_fd_sc_hd__clkbuf_2
X_4270_ _1894_ _1897_ VSS VSS VCC VCC _1898_ sky130_fd_sc_hd__nor2_1
X_3221_ _1166_ _1169_ VSS VSS VCC VCC _1170_ sky130_fd_sc_hd__nand2_2
X_3152_ _1109_ _1110_ VSS VSS VCC VCC net206 sky130_fd_sc_hd__nor2_8
X_3083_ _0798_ _0801_ _0788_ _0800_ net454 net629 VSS VSS VCC VCC _1045_ sky130_fd_sc_hd__mux4_1
X_3985_ u_wr_mux.i_reg_data2\[29\] net165 net391 VSS VSS VCC VCC _0147_ sky130_fd_sc_hd__mux2_1
X_2936_ net664 net667 net670 net673 net637 net625 VSS VSS VCC VCC _0906_ sky130_fd_sc_hd__mux4_1
X_2867_ net458 net650 VSS VSS VCC VCC _0839_ sky130_fd_sc_hd__and2_1
X_4606_ _1868_ _2163_ net473 _2166_ VSS VSS VCC VCC _2167_ sky130_fd_sc_hd__a31o_1
X_2798_ _0770_ _0771_ net622 VSS VSS VCC VCC _0772_ sky130_fd_sc_hd__mux2_1
X_4537_ u_muldiv.quotient_msk\[25\] net475 net332 u_muldiv.quotient_msk\[26\] vssd1
+ vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__a22o_1
X_4468_ u_muldiv.o_div\[21\] _2066_ u_muldiv.o_div\[22\] VSS VSS VCC VCC _2075_
+ sky130_fd_sc_hd__o21ai_1
X_3419_ net575 u_pc_sel.i_pc_next\[1\] _1314_ _1315_ VSS VSS VCC VCC net256
+ sky130_fd_sc_hd__a22o_2
X_4399_ u_muldiv.o_div\[7\] u_muldiv.o_div\[8\] _2012_ VSS VSS VCC VCC _2020_
+ sky130_fd_sc_hd__or3b_2
X_3770_ net139 net514 VSS VSS VCC VCC _1613_ sky130_fd_sc_hd__nand2b_1
X_2721_ net448 net594 VSS VSS VCC VCC _0696_ sky130_fd_sc_hd__nand2_1
X_2652_ _0609_ _0610_ _0613_ _0625_ _0615_ VSS VSS VCC VCC _0627_ sky130_fd_sc_hd__a32oi_4
Xclkbuf_4_2__f_i_clk clknet_2_0_0_i_clk VSS VSS VCC VCC clknet_4_2__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5371_ clknet_leaf_154_i_clk _0398_ VSS VSS VCC VCC u_muldiv.mul\[50\] sky130_fd_sc_hd__dfxtp_1
X_2583_ net447 net716 _0556_ VSS VSS VCC VCC _0558_ sky130_fd_sc_hd__a21oi_1
X_4322_ _1948_ _1949_ VSS VSS VCC VCC _1950_ sky130_fd_sc_hd__nand2_1
X_4253_ _1844_ _1876_ _1877_ _1880_ VSS VSS VCC VCC _1881_ sky130_fd_sc_hd__and4_1
X_3204_ op_cnt\[1\] op_cnt\[2\] op_cnt\[3\] VSS VSS VCC VCC _1159_ sky130_fd_sc_hd__and3_1
X_4184_ u_muldiv.mul\[14\] u_muldiv.mul\[13\] net404 VSS VSS VCC VCC _0228_
+ sky130_fd_sc_hd__mux2_1
X_3135_ _1076_ _1094_ net735 VSS VSS VCC VCC _1095_ sky130_fd_sc_hd__a21oi_4
X_3066_ _1026_ _1027_ VSS VSS VCC VCC _1029_ sky130_fd_sc_hd__nand2_2
X_3968_ u_wr_mux.i_reg_data2\[12\] net147 net389 VSS VSS VCC VCC _0130_ sky130_fd_sc_hd__mux2_1
X_2919_ _0889_ VSS VSS VCC VCC net199 sky130_fd_sc_hd__clkinv_8
X_3899_ u_bits.i_op2\[30\] u_bits.i_op2\[28\] net548 VSS VSS VCC VCC _1706_
+ sky130_fd_sc_hd__mux2_1
Xfanout620 net621 VSS VSS VCC VCC net620 sky130_fd_sc_hd__buf_4
Xfanout631 net633 VSS VSS VCC VCC net631 sky130_fd_sc_hd__clkbuf_4
Xfanout642 net644 VSS VSS VCC VCC net642 sky130_fd_sc_hd__clkbuf_8
Xfanout653 u_bits.i_op1\[30\] VSS VSS VCC VCC net653 sky130_fd_sc_hd__buf_6
Xfanout664 net666 VSS VSS VCC VCC net664 sky130_fd_sc_hd__buf_4
Xfanout675 u_bits.i_op1\[20\] VSS VSS VCC VCC net675 sky130_fd_sc_hd__buf_8
Xfanout686 net687 VSS VSS VCC VCC net686 sky130_fd_sc_hd__clkbuf_8
Xfanout697 net698 VSS VSS VCC VCC net697 sky130_fd_sc_hd__buf_4
X_4940_ _1167_ _1168_ net401 VSS VSS VCC VCC _0384_ sky130_fd_sc_hd__a21oi_1
X_4871_ u_muldiv.dividend\[29\] net316 _2408_ VSS VSS VCC VCC _0342_ sky130_fd_sc_hd__o21a_1
X_3822_ net596 net728 _1648_ _1647_ VSS VSS VCC VCC _0053_ sky130_fd_sc_hd__o22a_1
X_3753_ net678 net55 net391 VSS VSS VCC VCC _0022_ sky130_fd_sc_hd__mux2_1
X_2704_ _0674_ _0675_ _0677_ VSS VSS VCC VCC _0679_ sky130_fd_sc_hd__o21a_1
X_3684_ net561 _1562_ _1563_ net348 VSS VSS VCC VCC _1564_ sky130_fd_sc_hd__o211a_1
X_2635_ net518 net525 _0608_ VSS VSS VCC VCC _0610_ sky130_fd_sc_hd__o21ai_2
Xoutput201 net201 VSS VSS VCC VCC o_add[26] sky130_fd_sc_hd__buf_2
Xoutput212 net212 VSS VSS VCC VCC o_add[7] sky130_fd_sc_hd__buf_2
Xoutput223 net223 VSS VSS VCC VCC o_pc_target[13] sky130_fd_sc_hd__buf_2
X_5354_ clknet_leaf_103_i_clk _0381_ VSS VSS VCC VCC u_muldiv.mul\[33\] sky130_fd_sc_hd__dfxtp_1
Xoutput234 net234 VSS VSS VCC VCC o_pc_target[9] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VSS VSS VCC VCC o_result[0] sky130_fd_sc_hd__buf_2
X_2566_ net452 net537 _0460_ _0539_ VSS VSS VCC VCC _0541_ sky130_fd_sc_hd__o22ai_1
Xoutput256 net256 VSS VSS VCC VCC o_result[1] sky130_fd_sc_hd__buf_2
Xoutput267 net267 VSS VSS VCC VCC o_result[2] sky130_fd_sc_hd__buf_2
X_4305_ _1928_ _1930_ _1931_ VSS VSS VCC VCC _1933_ sky130_fd_sc_hd__and3_1
Xoutput278 net278 VSS VSS VCC VCC o_to_trap sky130_fd_sc_hd__buf_2
Xoutput289 net289 VSS VSS VCC VCC o_wdata[19] sky130_fd_sc_hd__buf_2
X_5285_ clknet_leaf_7_i_clk _0313_ VSS VSS VCC VCC u_muldiv.quotient_msk\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_2497_ _0471_ _0468_ VSS VSS VCC VCC _0472_ sky130_fd_sc_hd__nand2_1
X_4236_ u_muldiv.divisor\[3\] _0441_ _1863_ VSS VSS VCC VCC _1864_ sky130_fd_sc_hd__o21a_1
X_4167_ net549 net499 net203 VSS VSS VCC VCC _0211_ sky130_fd_sc_hd__o21a_1
X_3118_ net612 _1077_ net347 VSS VSS VCC VCC _1078_ sky130_fd_sc_hd__o21a_1
X_4098_ u_bits.i_op2\[22\] _1803_ _1804_ VSS VSS VCC VCC _1805_ sky130_fd_sc_hd__o21ba_1
X_3049_ net623 _0859_ _1012_ VSS VSS VCC VCC _1013_ sky130_fd_sc_hd__o21ai_2
Xfanout450 net451 VSS VSS VCC VCC net450 sky130_fd_sc_hd__buf_4
Xfanout461 u_bits.i_op1\[0\] VSS VSS VCC VCC net461 sky130_fd_sc_hd__buf_2
Xfanout472 net474 VSS VSS VCC VCC net472 sky130_fd_sc_hd__clkbuf_4
Xfanout483 net487 VSS VSS VCC VCC net483 sky130_fd_sc_hd__buf_4
Xfanout494 net495 VSS VSS VCC VCC net494 sky130_fd_sc_hd__clkbuf_4
X_5070_ clknet_leaf_173_i_clk _0103_ VSS VSS VCC VCC net220 sky130_fd_sc_hd__dfxtp_1
X_4021_ net599 _1742_ _1743_ VSS VSS VCC VCC _1744_ sky130_fd_sc_hd__o21ba_1
X_4923_ u_muldiv.divisor\[30\] net477 net333 u_muldiv.divisor\[31\] vssd1 vssd1 vccd1
+ vccd1 _0375_ sky130_fd_sc_hd__a22o_1
X_4854_ _2389_ _2390_ _2392_ VSS VSS VCC VCC _2393_ sky130_fd_sc_hd__o21ai_1
X_3805_ net504 net104 net720 VSS VSS VCC VCC _1636_ sky130_fd_sc_hd__a21o_1
X_4785_ net670 _2329_ VSS VSS VCC VCC _2330_ sky130_fd_sc_hd__nor2_1
X_3736_ u_bits.i_op1\[2\] net67 net389 VSS VSS VCC VCC _0005_ sky130_fd_sc_hd__mux2_1
X_3667_ net628 net346 _0847_ net605 VSS VSS VCC VCC _1548_ sky130_fd_sc_hd__o31a_1
X_2618_ _0591_ _0592_ VSS VSS VCC VCC _0593_ sky130_fd_sc_hd__nand2_1
X_3598_ _1047_ net345 net412 _1483_ _1480_ VSS VSS VCC VCC _1484_ sky130_fd_sc_hd__a2111oi_1
X_5337_ clknet_leaf_163_i_clk _0365_ VSS VSS VCC VCC u_muldiv.divisor\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_2549_ net685 u_muldiv.add_prev\[16\] net536 VSS VSS VCC VCC _0524_ sky130_fd_sc_hd__mux2_1
X_5268_ clknet_leaf_128_i_clk _0296_ VSS VSS VCC VCC u_muldiv.quotient_msk\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_4219_ u_muldiv.divisor\[5\] u_muldiv.dividend\[5\] VSS VSS VCC VCC _1847_
+ sky130_fd_sc_hd__and2b_1
X_5199_ clknet_leaf_154_i_clk _0231_ VSS VSS VCC VCC u_muldiv.mul\[16\] sky130_fd_sc_hd__dfxtp_1
X_4570_ net497 _2132_ _2133_ _1720_ VSS VSS VCC VCC _2134_ sky130_fd_sc_hd__o31a_1
X_3521_ _1410_ _1411_ _0838_ _0842_ net616 net609 VSS VSS VCC VCC _1412_ sky130_fd_sc_hd__mux4_2
X_3452_ net452 net568 net712 VSS VSS VCC VCC _1347_ sky130_fd_sc_hd__or3b_1
X_3383_ net565 _0846_ net350 VSS VSS VCC VCC _1281_ sky130_fd_sc_hd__o21a_1
X_5122_ clknet_leaf_16_i_clk _0154_ VSS VSS VCC VCC u_muldiv.divisor\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_5053_ clknet_leaf_163_i_clk _0086_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4004_ u_muldiv.divisor\[33\] net478 net333 u_muldiv.divisor\[34\] _1730_ vssd1 vssd1
+ vccd1 vccd1 _0153_ sky130_fd_sc_hd__a221o_1
X_4906_ u_muldiv.divisor\[13\] net490 net338 u_muldiv.divisor\[14\] vssd1 vssd1 vccd1
+ vccd1 _0358_ sky130_fd_sc_hd__a22o_1
X_4837_ _1953_ _2376_ net465 VSS VSS VCC VCC _2377_ sky130_fd_sc_hd__o21ai_1
X_4768_ _1937_ _1939_ _2313_ VSS VSS VCC VCC _2314_ sky130_fd_sc_hd__or3_1
X_3719_ u_muldiv.mul\[53\] net361 net357 u_muldiv.mul\[21\] _1595_ vssd1 vssd1 vccd1
+ vccd1 _1596_ sky130_fd_sc_hd__a221o_2
X_4699_ u_muldiv.dividend\[14\] net326 net377 _2251_ VSS VSS VCC VCC _0327_
+ sky130_fd_sc_hd__a31o_1
X_2952_ net445 u_bits.i_op2\[25\] _0464_ net663 VSS VSS VCC VCC _0921_ sky130_fd_sc_hd__a22o_1
X_2883_ net456 _0852_ _0854_ VSS VSS VCC VCC _0855_ sky130_fd_sc_hd__o21ai_1
X_4622_ u_muldiv.dividend\[7\] _2161_ u_muldiv.dividend\[8\] VSS VSS VCC VCC
+ _2181_ sky130_fd_sc_hd__o21ai_1
X_4553_ net464 _1992_ _2118_ VSS VSS VCC VCC _0314_ sky130_fd_sc_hd__a21o_1
X_3504_ _0905_ _1316_ _1318_ _0908_ VSS VSS VCC VCC _1396_ sky130_fd_sc_hd__o22a_1
X_4484_ net315 _2085_ _2087_ VSS VSS VCC VCC _0276_ sky130_fd_sc_hd__a21oi_1
X_3435_ _0422_ _1329_ _1330_ net354 net205 VSS VSS VCC VCC _1331_ sky130_fd_sc_hd__a32o_1
X_3366_ net417 net183 net568 net194 VSS VSS VCC VCC net313 sky130_fd_sc_hd__o2bb2a_4
X_5105_ clknet_leaf_60_i_clk _0138_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_3297_ _1217_ _1226_ VSS VSS VCC VCC _1227_ sky130_fd_sc_hd__nor2_1
X_5036_ clknet_leaf_26_i_clk _0069_ VSS VSS VCC VCC u_bits.i_op2\[25\] sky130_fd_sc_hd__dfxtp_2
Xinput101 i_op2[31] VSS VSS VCC VCC net101 sky130_fd_sc_hd__clkbuf_1
Xinput112 i_pc_next[13] VSS VSS VCC VCC net112 sky130_fd_sc_hd__clkbuf_1
Xinput123 i_pc_next[9] VSS VSS VCC VCC net123 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput134 i_pc_target[5] VSS VSS VCC VCC net134 sky130_fd_sc_hd__clkbuf_4
Xinput145 i_reg_data2[10] VSS VSS VCC VCC net145 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput156 i_reg_data2[20] VSS VSS VCC VCC net156 sky130_fd_sc_hd__clkbuf_1
Xinput167 i_reg_data2[30] VSS VSS VCC VCC net167 sky130_fd_sc_hd__clkbuf_2
Xinput178 i_res_src[1] VSS VSS VCC VCC net178 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_132_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_132_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3220_ _0591_ _0592_ _0584_ VSS VSS VCC VCC _1169_ sky130_fd_sc_hd__a21o_1
X_3151_ _1030_ _1069_ _1035_ _1108_ _1100_ VSS VSS VCC VCC _1110_ sky130_fd_sc_hd__o311a_2
X_3082_ net457 _0898_ _1043_ VSS VSS VCC VCC _1044_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_leaf_147_i_clk clknet_4_8__leaf_i_clk VSS VSS VCC VCC clknet_leaf_147_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3984_ u_wr_mux.i_reg_data2\[28\] net164 net398 VSS VSS VCC VCC _0146_ sky130_fd_sc_hd__mux2_1
X_2935_ net452 net623 VSS VSS VCC VCC _0905_ sky130_fd_sc_hd__nand2_8
X_2866_ _0836_ _0837_ net456 VSS VSS VCC VCC _0838_ sky130_fd_sc_hd__mux2_1
X_4605_ net707 _2164_ _2165_ VSS VSS VCC VCC _2166_ sky130_fd_sc_hd__o21a_1
X_2797_ net660 net658 net657 net655 net639 net625 VSS VSS VCC VCC _0771_ sky130_fd_sc_hd__mux4_1
X_4536_ u_muldiv.quotient_msk\[24\] net475 net332 u_muldiv.quotient_msk\[25\] vssd1
+ vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__a22o_1
X_4467_ u_muldiv.o_div\[19\] _2059_ _2073_ _0456_ VSS VSS VCC VCC _2074_ sky130_fd_sc_hd__nand4b_4
X_3418_ net17 net729 net575 VSS VSS VCC VCC _1315_ sky130_fd_sc_hd__o21ba_1
X_4398_ u_muldiv.o_div\[5\] u_muldiv.o_div\[6\] u_muldiv.o_div\[7\] _2006_ vssd1 vssd1
+ vccd1 vccd1 _2019_ sky130_fd_sc_hd__nor4_1
X_3349_ u_wr_mux.i_reg_data2\[8\] _0764_ _1258_ VSS VSS VCC VCC net295 sky130_fd_sc_hd__a21o_4
X_5019_ clknet_leaf_55_i_clk _0052_ VSS VSS VCC VCC u_bits.i_op2\[8\] sky130_fd_sc_hd__dfxtp_4
X_2720_ _0693_ _0694_ VSS VSS VCC VCC _0695_ sky130_fd_sc_hd__and2_1
X_2651_ _0622_ _0623_ _0618_ _0619_ VSS VSS VCC VCC _0626_ sky130_fd_sc_hd__o211ai_2
Xclkbuf_leaf_17_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_17_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2582_ net447 net716 VSS VSS VCC VCC _0557_ sky130_fd_sc_hd__and2_1
X_5370_ clknet_leaf_107_i_clk _0397_ VSS VSS VCC VCC u_muldiv.mul\[49\] sky130_fd_sc_hd__dfxtp_1
X_4321_ u_muldiv.dividend\[26\] u_muldiv.divisor\[26\] VSS VSS VCC VCC _1949_
+ sky130_fd_sc_hd__nand2b_1
X_4252_ u_muldiv.divisor\[9\] u_muldiv.dividend\[9\] VSS VSS VCC VCC _1880_
+ sky130_fd_sc_hd__nand2b_1
X_3203_ op_cnt\[1\] _1157_ net548 VSS VSS VCC VCC _1158_ sky130_fd_sc_hd__or3b_1
X_4183_ u_muldiv.mul\[13\] u_muldiv.mul\[12\] net403 VSS VSS VCC VCC _0227_
+ sky130_fd_sc_hd__mux2_1
X_3134_ _1093_ _1092_ net204 net355 net527 VSS VSS VCC VCC _1094_ sky130_fd_sc_hd__a221o_1
X_3065_ _1027_ _1026_ VSS VSS VCC VCC _1028_ sky130_fd_sc_hd__or2_1
X_3967_ u_wr_mux.i_reg_data2\[11\] net146 net386 VSS VSS VCC VCC _0129_ sky130_fd_sc_hd__mux2_1
X_2918_ _0877_ _0887_ VSS VSS VCC VCC _0889_ sky130_fd_sc_hd__xor2_4
X_3898_ u_bits.i_op2\[28\] net727 _1705_ _1704_ VSS VSS VCC VCC _0072_ sky130_fd_sc_hd__o22a_1
X_2849_ net669 u_muldiv.add_prev\[23\] net533 VSS VSS VCC VCC _0822_ sky130_fd_sc_hd__mux2_1
X_4519_ u_muldiv.quotient_msk\[7\] net493 net339 u_muldiv.quotient_msk\[8\] vssd1
+ vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__a22o_1
Xfanout610 u_bits.i_op2\[4\] VSS VSS VCC VCC net610 sky130_fd_sc_hd__clkbuf_4
Xfanout621 net622 VSS VSS VCC VCC net621 sky130_fd_sc_hd__buf_4
Xfanout632 net633 VSS VSS VCC VCC net632 sky130_fd_sc_hd__buf_4
Xfanout643 net644 VSS VSS VCC VCC net643 sky130_fd_sc_hd__buf_4
Xfanout654 u_bits.i_op1\[29\] VSS VSS VCC VCC net654 sky130_fd_sc_hd__buf_6
Xfanout665 net666 VSS VSS VCC VCC net665 sky130_fd_sc_hd__clkbuf_2
Xfanout676 u_bits.i_op1\[20\] VSS VSS VCC VCC net676 sky130_fd_sc_hd__clkbuf_4
Xfanout687 u_bits.i_op1\[15\] VSS VSS VCC VCC net687 sky130_fd_sc_hd__buf_8
Xfanout698 u_bits.i_op1\[10\] VSS VSS VCC VCC net698 sky130_fd_sc_hd__buf_6
X_4870_ _2399_ _2400_ _2407_ net316 VSS VSS VCC VCC _2408_ sky130_fd_sc_hd__o211ai_1
X_3821_ net512 net108 net721 VSS VSS VCC VCC _1648_ sky130_fd_sc_hd__a21o_1
X_3752_ net680 net54 net386 VSS VSS VCC VCC _0021_ sky130_fd_sc_hd__mux2_1
X_2703_ _0677_ VSS VSS VCC VCC _0678_ sky130_fd_sc_hd__inv_2
X_3683_ net588 net680 VSS VSS VCC VCC _1563_ sky130_fd_sc_hd__or2_1
X_2634_ net540 _0426_ net431 _0607_ VSS VSS VCC VCC _0609_ sky130_fd_sc_hd__o211ai_4
Xoutput202 net202 VSS VSS VCC VCC o_add[27] sky130_fd_sc_hd__buf_2
Xoutput213 net213 VSS VSS VCC VCC o_add[8] sky130_fd_sc_hd__buf_2
Xoutput224 net224 VSS VSS VCC VCC o_pc_target[14] sky130_fd_sc_hd__buf_2
Xoutput235 net235 VSS VSS VCC VCC o_rd[0] sky130_fd_sc_hd__buf_2
X_2565_ net647 net551 _0538_ net423 VSS VSS VCC VCC _0540_ sky130_fd_sc_hd__o211ai_2
X_5353_ clknet_leaf_104_i_clk _0380_ VSS VSS VCC VCC u_muldiv.mul\[32\] sky130_fd_sc_hd__dfxtp_1
Xoutput246 net246 VSS VSS VCC VCC o_result[10] sky130_fd_sc_hd__buf_2
Xoutput257 net257 VSS VSS VCC VCC o_result[20] sky130_fd_sc_hd__buf_2
X_4304_ _1930_ _1931_ VSS VSS VCC VCC _1932_ sky130_fd_sc_hd__and2_1
Xoutput268 net268 VSS VSS VCC VCC o_result[30] sky130_fd_sc_hd__buf_2
Xoutput279 net279 VSS VSS VCC VCC o_wdata[0] sky130_fd_sc_hd__buf_2
X_2496_ _0466_ net430 _0465_ _0469_ VSS VSS VCC VCC _0471_ sky130_fd_sc_hd__o31a_1
X_5284_ clknet_leaf_7_i_clk _0312_ VSS VSS VCC VCC u_muldiv.quotient_msk\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_4235_ _0417_ net463 _1853_ _1861_ VSS VSS VCC VCC _1863_ sky130_fd_sc_hd__o211ai_2
X_4166_ _1000_ _1001_ net400 VSS VSS VCC VCC _0210_ sky130_fd_sc_hd__and3_1
X_3117_ net619 _0931_ _0773_ VSS VSS VCC VCC _1077_ sky130_fd_sc_hd__o21a_1
X_4097_ u_bits.i_op2\[22\] _1803_ net484 net468 VSS VSS VCC VCC _1804_ sky130_fd_sc_hd__a211o_1
X_3048_ net456 _0853_ VSS VSS VCC VCC _1012_ sky130_fd_sc_hd__or2_1
X_4999_ clknet_leaf_148_i_clk _0032_ VSS VSS VCC VCC u_bits.i_op1\[29\] sky130_fd_sc_hd__dfxtp_4
Xfanout440 _0434_ VSS VSS VCC VCC net440 sky130_fd_sc_hd__buf_6
Xfanout451 _0421_ VSS VSS VCC VCC net451 sky130_fd_sc_hd__clkbuf_8
Xfanout462 u_muldiv.dividend\[17\] VSS VSS VCC VCC net462 sky130_fd_sc_hd__buf_4
Xfanout473 net474 VSS VSS VCC VCC net473 sky130_fd_sc_hd__buf_4
Xfanout484 net486 VSS VSS VCC VCC net484 sky130_fd_sc_hd__clkbuf_4
Xfanout495 u_muldiv.i_on_end VSS VSS VCC VCC net495 sky130_fd_sc_hd__clkbuf_4
X_4020_ _1741_ net379 net599 net329 VSS VSS VCC VCC _1743_ sky130_fd_sc_hd__a31o_1
X_4922_ u_muldiv.divisor\[29\] net478 net333 u_muldiv.divisor\[30\] vssd1 vssd1 vccd1
+ vccd1 _0374_ sky130_fd_sc_hd__a22o_1
X_4853_ _1960_ _1966_ _2391_ VSS VSS VCC VCC _2392_ sky130_fd_sc_hd__a21o_1
X_3804_ net504 _1634_ VSS VSS VCC VCC _1635_ sky130_fd_sc_hd__and2b_1
X_4784_ net672 _2316_ net371 VSS VSS VCC VCC _2329_ sky130_fd_sc_hd__o21a_1
X_3735_ u_bits.i_op1\[1\] net56 net390 VSS VSS VCC VCC _0004_ sky130_fd_sc_hd__mux2_1
X_3666_ net604 _1296_ net327 VSS VSS VCC VCC _1547_ sky130_fd_sc_hd__o21ai_1
X_2617_ _0586_ _0588_ _0590_ _0587_ VSS VSS VCC VCC _0592_ sky130_fd_sc_hd__a211o_1
X_3597_ net593 net693 _1482_ VSS VSS VCC VCC _1483_ sky130_fd_sc_hd__o21a_1
X_5336_ clknet_leaf_163_i_clk _0364_ VSS VSS VCC VCC u_muldiv.divisor\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_2548_ _0521_ net432 VSS VSS VCC VCC _0523_ sky130_fd_sc_hd__nand2_1
X_5267_ clknet_leaf_128_i_clk _0295_ VSS VSS VCC VCC u_muldiv.quotient_msk\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_2479_ u_muldiv.o_div\[12\] VSS VSS VCC VCC _0454_ sky130_fd_sc_hd__inv_2
X_4218_ u_muldiv.divisor\[7\] u_muldiv.dividend\[7\] VSS VSS VCC VCC _1846_
+ sky130_fd_sc_hd__nand2b_1
X_5198_ clknet_leaf_155_i_clk _0230_ VSS VSS VCC VCC u_muldiv.mul\[15\] sky130_fd_sc_hd__dfxtp_1
X_4149_ _1185_ _1189_ net402 VSS VSS VCC VCC _0193_ sky130_fd_sc_hd__and3_1
X_3520_ _1337_ _1339_ net457 VSS VSS VCC VCC _1411_ sky130_fd_sc_hd__mux2_1
X_3451_ net609 _1338_ _1345_ VSS VSS VCC VCC _1346_ sky130_fd_sc_hd__a21o_1
X_3382_ net628 net620 net613 _0791_ VSS VSS VCC VCC _1280_ sky130_fd_sc_hd__or4_1
X_5121_ clknet_leaf_16_i_clk _0153_ VSS VSS VCC VCC u_muldiv.divisor\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_5052_ clknet_leaf_137_i_clk _0085_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_4003_ net624 _1728_ _1729_ VSS VSS VCC VCC _1730_ sky130_fd_sc_hd__o21ba_1
X_4905_ u_muldiv.divisor\[12\] net490 net338 u_muldiv.divisor\[13\] vssd1 vssd1 vccd1
+ vccd1 _0357_ sky130_fd_sc_hd__a22o_1
X_4836_ _1948_ _2367_ VSS VSS VCC VCC _2376_ sky130_fd_sc_hd__nand2_1
X_4767_ _1936_ _1925_ _1934_ VSS VSS VCC VCC _2313_ sky130_fd_sc_hd__o21bai_1
X_3718_ u_muldiv.dividend\[21\] net419 net364 u_muldiv.o_div\[21\] net442 vssd1 vssd1
+ vccd1 vccd1 _1595_ sky130_fd_sc_hd__a221o_1
X_4698_ _2250_ net437 net326 net377 _2244_ VSS VSS VCC VCC _2251_ sky130_fd_sc_hd__a221oi_1
X_3649_ net12 net730 net576 VSS VSS VCC VCC _1532_ sky130_fd_sc_hd__o21ba_1
X_5319_ clknet_leaf_91_i_clk _0347_ VSS VSS VCC VCC u_muldiv.divisor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_3_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_3_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_2951_ _0876_ _0887_ _0875_ VSS VSS VCC VCC _0920_ sky130_fd_sc_hd__o21ai_2
X_2882_ net623 _0853_ VSS VSS VCC VCC _0854_ sky130_fd_sc_hd__or2_1
X_4621_ u_muldiv.dividend\[7\] u_muldiv.dividend\[8\] _2161_ VSS VSS VCC VCC
+ _2180_ sky130_fd_sc_hd__or3_2
X_4552_ net498 _2109_ _2112_ _2117_ net322 VSS VSS VCC VCC _2118_ sky130_fd_sc_hd__a221oi_1
X_3503_ net622 _1317_ _1394_ VSS VSS VCC VCC _1395_ sky130_fd_sc_hd__o21ai_1
X_4483_ net315 _2086_ u_muldiv.o_div\[25\] VSS VSS VCC VCC _2087_ sky130_fd_sc_hd__a21oi_1
X_3434_ net621 net715 _0781_ net441 VSS VSS VCC VCC _1330_ sky130_fd_sc_hd__a211o_1
X_3365_ net183 _0758_ net560 _1213_ VSS VSS VCC VCC net312 sky130_fd_sc_hd__o22a_2
X_5104_ clknet_leaf_72_i_clk _0137_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[19\]
+ sky130_fd_sc_hd__dfxtp_4
X_3296_ _1181_ _1190_ _1198_ _1219_ VSS VSS VCC VCC _1226_ sky130_fd_sc_hd__nand4_1
X_5035_ clknet_leaf_31_i_clk _0068_ VSS VSS VCC VCC u_bits.i_op2\[24\] sky130_fd_sc_hd__dfxtp_4
X_4819_ net476 _2359_ _2360_ _1720_ VSS VSS VCC VCC _2361_ sky130_fd_sc_hd__o31a_1
Xinput102 i_op2[3] VSS VSS VCC VCC net102 sky130_fd_sc_hd__clkbuf_2
Xinput113 i_pc_next[14] VSS VSS VCC VCC net113 sky130_fd_sc_hd__clkbuf_1
Xinput124 i_pc_target[10] VSS VSS VCC VCC net124 sky130_fd_sc_hd__buf_4
Xinput135 i_pc_target[6] VSS VSS VCC VCC net135 sky130_fd_sc_hd__buf_6
Xinput146 i_reg_data2[11] VSS VSS VCC VCC net146 sky130_fd_sc_hd__clkbuf_1
Xinput157 i_reg_data2[21] VSS VSS VCC VCC net157 sky130_fd_sc_hd__clkbuf_1
Xinput168 i_reg_data2[31] VSS VSS VCC VCC net168 sky130_fd_sc_hd__clkbuf_1
Xinput179 i_res_src[2] VSS VSS VCC VCC net179 sky130_fd_sc_hd__buf_4
X_3150_ _1099_ _1100_ _1108_ VSS VSS VCC VCC _1109_ sky130_fd_sc_hd__a21oi_4
X_3081_ net623 net460 _0840_ VSS VSS VCC VCC _1043_ sky130_fd_sc_hd__and3_1
X_3983_ u_wr_mux.i_reg_data2\[27\] net163 net391 VSS VSS VCC VCC _0145_ sky130_fd_sc_hd__mux2_1
X_2934_ net675 net677 net679 net682 net642 net627 VSS VSS VCC VCC _0904_ sky130_fd_sc_hd__mux4_2
X_2865_ net669 net666 net663 net661 net641 net636 VSS VSS VCC VCC _0837_ sky130_fd_sc_hd__mux4_2
X_4604_ net707 _2164_ net473 VSS VSS VCC VCC _2165_ sky130_fd_sc_hd__a21oi_1
X_2796_ net671 net668 net665 net663 net639 net625 VSS VSS VCC VCC _0770_ sky130_fd_sc_hd__mux4_1
X_4535_ u_muldiv.quotient_msk\[23\] net480 net334 u_muldiv.quotient_msk\[24\] vssd1
+ vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__a22o_1
X_4466_ u_muldiv.o_div\[22\] u_muldiv.o_div\[21\] VSS VSS VCC VCC _2073_ sky130_fd_sc_hd__nor2_1
X_3417_ _1308_ _1310_ _1313_ net733 VSS VSS VCC VCC _1314_ sky130_fd_sc_hd__a211o_4
X_4397_ net322 _2016_ _2018_ VSS VSS VCC VCC _0258_ sky130_fd_sc_hd__o21a_1
X_3348_ net563 u_wr_mux.i_reg_data2\[24\] net416 net279 VSS VSS VCC VCC _1258_
+ sky130_fd_sc_hd__a22o_1
X_3279_ _0568_ _0569_ VSS VSS VCC VCC _1212_ sky130_fd_sc_hd__nand2_2
X_5018_ clknet_leaf_27_i_clk _0051_ VSS VSS VCC VCC u_bits.i_op2\[7\] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0_i_clk i_clk VSS VSS VCC VCC clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_2650_ _0622_ _0623_ _0618_ _0619_ VSS VSS VCC VCC _0625_ sky130_fd_sc_hd__o211a_2
X_2581_ net538 u_muldiv.add_prev\[2\] VSS VSS VCC VCC _0556_ sky130_fd_sc_hd__and2_1
X_4320_ u_muldiv.divisor\[26\] u_muldiv.dividend\[26\] VSS VSS VCC VCC _1948_
+ sky130_fd_sc_hd__nand2b_1
X_4251_ _1875_ _1878_ VSS VSS VCC VCC _1879_ sky130_fd_sc_hd__or2_1
X_3202_ op_cnt\[2\] op_cnt\[3\] op_cnt\[4\] op_cnt\[5\] VSS VSS VCC VCC _1157_
+ sky130_fd_sc_hd__or4b_1
X_4182_ u_muldiv.mul\[12\] u_muldiv.mul\[11\] net403 VSS VSS VCC VCC _0226_
+ sky130_fd_sc_hd__mux2_1
X_3133_ net410 _1083_ net522 VSS VSS VCC VCC _1093_ sky130_fd_sc_hd__a21oi_1
X_3064_ net657 u_muldiv.add_prev\[28\] net533 VSS VSS VCC VCC _1027_ sky130_fd_sc_hd__mux2_1
X_3966_ u_wr_mux.i_reg_data2\[10\] net145 net392 VSS VSS VCC VCC _0128_ sky130_fd_sc_hd__mux2_1
X_2917_ _0880_ _0743_ _0885_ VSS VSS VCC VCC _0888_ sky130_fd_sc_hd__o21ai_2
X_3897_ net509 net97 net721 VSS VSS VCC VCC _1705_ sky130_fd_sc_hd__a21o_1
X_2848_ net732 net20 _0821_ VSS VSS VCC VCC net259 sky130_fd_sc_hd__o21a_2
X_2779_ _0753_ VSS VSS VCC VCC net197 sky130_fd_sc_hd__inv_2
X_4518_ u_muldiv.quotient_msk\[6\] net493 net342 u_muldiv.quotient_msk\[7\] vssd1
+ vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__a22o_1
X_4449_ u_muldiv.o_div\[16\] u_muldiv.o_div\[17\] u_muldiv.o_div\[18\] _2050_ net490
+ VSS VSS VCC VCC _2060_ sky130_fd_sc_hd__o41a_1
Xfanout600 u_bits.i_op2\[5\] VSS VSS VCC VCC net600 sky130_fd_sc_hd__buf_6
Xfanout611 net612 VSS VSS VCC VCC net611 sky130_fd_sc_hd__buf_4
Xfanout622 u_bits.i_op2\[2\] VSS VSS VCC VCC net622 sky130_fd_sc_hd__buf_2
Xfanout633 u_bits.i_op2\[1\] VSS VSS VCC VCC net633 sky130_fd_sc_hd__buf_4
Xfanout644 net645 VSS VSS VCC VCC net644 sky130_fd_sc_hd__buf_6
Xfanout655 u_bits.i_op1\[29\] VSS VSS VCC VCC net655 sky130_fd_sc_hd__buf_4
Xfanout666 u_bits.i_op1\[24\] VSS VSS VCC VCC net666 sky130_fd_sc_hd__buf_6
Xfanout677 u_bits.i_op1\[19\] VSS VSS VCC VCC net677 sky130_fd_sc_hd__buf_4
Xfanout688 net689 VSS VSS VCC VCC net688 sky130_fd_sc_hd__buf_4
Xfanout699 net700 VSS VSS VCC VCC net699 sky130_fd_sc_hd__buf_4
X_3820_ net513 _1646_ VSS VSS VCC VCC _1647_ sky130_fd_sc_hd__and2b_1
X_3751_ net682 net53 net386 VSS VSS VCC VCC _0020_ sky130_fd_sc_hd__mux2_1
X_2702_ net689 u_muldiv.add_prev\[14\] net542 VSS VSS VCC VCC _0677_ sky130_fd_sc_hd__mux2_2
X_3682_ net588 net680 VSS VSS VCC VCC _1562_ sky130_fd_sc_hd__nand2_1
X_2633_ net540 _0426_ _0607_ VSS VSS VCC VCC _0608_ sky130_fd_sc_hd__o21ai_1
Xoutput203 net203 VSS VSS VCC VCC o_add[28] sky130_fd_sc_hd__buf_2
Xoutput214 net214 VSS VSS VCC VCC o_add[9] sky130_fd_sc_hd__buf_2
X_5352_ clknet_4_12__leaf_i_clk _0379_ VSS VSS VCC VCC u_muldiv.mul\[31\]
+ sky130_fd_sc_hd__dfxtp_2
X_2564_ net646 net551 net714 net538 VSS VSS VCC VCC _0539_ sky130_fd_sc_hd__o211ai_2
Xoutput225 net225 VSS VSS VCC VCC o_pc_target[15] sky130_fd_sc_hd__buf_2
Xoutput236 net236 VSS VSS VCC VCC o_rd[1] sky130_fd_sc_hd__buf_2
Xoutput247 net247 VSS VSS VCC VCC o_result[11] sky130_fd_sc_hd__buf_2
Xoutput258 net258 VSS VSS VCC VCC o_result[21] sky130_fd_sc_hd__buf_2
X_4303_ u_muldiv.dividend\[23\] u_muldiv.divisor\[23\] VSS VSS VCC VCC _1931_
+ sky130_fd_sc_hd__nand2b_1
Xoutput269 net269 VSS VSS VCC VCC o_result[31] sky130_fd_sc_hd__buf_2
X_5283_ clknet_leaf_1_i_clk _0311_ VSS VSS VCC VCC u_muldiv.quotient_msk\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_2495_ _0467_ _0468_ _0469_ VSS VSS VCC VCC _0470_ sky130_fd_sc_hd__a21o_1
X_4234_ _0417_ net463 _1861_ VSS VSS VCC VCC _1862_ sky130_fd_sc_hd__o21a_1
X_4165_ net550 net500 net201 VSS VSS VCC VCC _0209_ sky130_fd_sc_hd__o21a_1
X_3116_ u_muldiv.mul\[61\] net440 _0758_ _1075_ VSS VSS VCC VCC _1076_ sky130_fd_sc_hd__a31o_1
X_4096_ u_bits.i_op2\[20\] u_bits.i_op2\[21\] _1795_ net380 VSS VSS VCC VCC
+ _1803_ sky130_fd_sc_hd__o31a_1
X_3047_ net457 net616 _0848_ _1010_ VSS VSS VCC VCC _1011_ sky130_fd_sc_hd__a31o_2
X_4998_ clknet_leaf_51_i_clk _0031_ VSS VSS VCC VCC u_bits.i_op1\[28\] sky130_fd_sc_hd__dfxtp_1
X_3949_ net550 net1 net389 VSS VSS VCC VCC _0112_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_78_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_78_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout430 _0458_ VSS VSS VCC VCC net430 sky130_fd_sc_hd__buf_4
Xfanout441 _0434_ VSS VSS VCC VCC net441 sky130_fd_sc_hd__buf_6
Xfanout452 _0421_ VSS VSS VCC VCC net452 sky130_fd_sc_hd__buf_6
Xfanout463 u_muldiv.dividend\[2\] VSS VSS VCC VCC net463 sky130_fd_sc_hd__buf_4
Xfanout474 u_muldiv.on_wait VSS VSS VCC VCC net474 sky130_fd_sc_hd__clkbuf_4
Xfanout485 net486 VSS VSS VCC VCC net485 sky130_fd_sc_hd__clkbuf_2
Xfanout496 net497 VSS VSS VCC VCC net496 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_16_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_16_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4921_ u_muldiv.divisor\[28\] net475 net332 u_muldiv.divisor\[29\] vssd1 vssd1 vccd1
+ vccd1 _0373_ sky130_fd_sc_hd__a22o_1
X_4852_ _1966_ _1960_ net465 VSS VSS VCC VCC _2391_ sky130_fd_sc_hd__o21ai_1
X_3803_ net599 net603 net546 VSS VSS VCC VCC _1634_ sky130_fd_sc_hd__mux2_1
X_4783_ _1928_ _2326_ _2327_ VSS VSS VCC VCC _2328_ sky130_fd_sc_hd__a21o_1
X_3734_ net39 net180 net512 VSS VSS VCC VCC _1610_ sky130_fd_sc_hd__and3b_4
X_3665_ u_muldiv.mul\[49\] net361 net360 u_muldiv.mul\[17\] VSS VSS VCC VCC
+ _1546_ sky130_fd_sc_hd__a22oi_1
X_2616_ _0587_ _0589_ _0590_ VSS VSS VCC VCC _0591_ sky130_fd_sc_hd__o21ai_4
X_3596_ net564 _1481_ net350 VSS VSS VCC VCC _1482_ sky130_fd_sc_hd__o21a_1
X_5335_ clknet_leaf_148_i_clk _0363_ VSS VSS VCC VCC u_muldiv.divisor\[18\]
+ sky130_fd_sc_hd__dfxtp_2
X_2547_ net536 _0428_ net517 net524 _0520_ VSS VSS VCC VCC _0522_ sky130_fd_sc_hd__o221ai_4
X_5266_ clknet_leaf_120_i_clk _0294_ VSS VSS VCC VCC u_muldiv.quotient_msk\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2478_ u_muldiv.o_div\[9\] VSS VSS VCC VCC _0453_ sky130_fd_sc_hd__inv_2
X_4217_ u_muldiv.dividend\[7\] u_muldiv.divisor\[7\] VSS VSS VCC VCC _1845_
+ sky130_fd_sc_hd__nand2b_1
X_5197_ clknet_leaf_107_i_clk _0229_ VSS VSS VCC VCC u_muldiv.mul\[14\] sky130_fd_sc_hd__dfxtp_1
X_4148_ _1179_ _1180_ net402 VSS VSS VCC VCC _0192_ sky130_fd_sc_hd__and3_1
X_4079_ _1788_ _1789_ VSS VSS VCC VCC _1790_ sky130_fd_sc_hd__nor2_1
X_3450_ net346 _1342_ net452 _1341_ _1344_ VSS VSS VCC VCC _1345_ sky130_fd_sc_hd__o221a_1
X_3381_ net640 net636 net624 net618 VSS VSS VCC VCC _1279_ sky130_fd_sc_hd__or4_1
X_5120_ clknet_leaf_16_i_clk _0152_ VSS VSS VCC VCC u_muldiv.divisor\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_5051_ clknet_4_0__leaf_i_clk _0084_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[9\]
+ sky130_fd_sc_hd__dfxtp_4
X_4002_ net624 _1728_ net478 net467 VSS VSS VCC VCC _1729_ sky130_fd_sc_hd__a211o_1
X_4904_ u_muldiv.divisor\[11\] net490 net338 u_muldiv.divisor\[12\] vssd1 vssd1 vccd1
+ vccd1 _0356_ sky130_fd_sc_hd__a22o_1
X_4835_ _2375_ u_muldiv.dividend\[26\] net323 VSS VSS VCC VCC _0339_ sky130_fd_sc_hd__mux2_1
X_4766_ u_muldiv.dividend\[20\] _1990_ _1991_ _2312_ VSS VSS VCC VCC _0333_
+ sky130_fd_sc_hd__a31o_1
X_3717_ net729 net18 _1594_ VSS VSS VCC VCC net257 sky130_fd_sc_hd__o21a_4
X_4697_ net469 _2248_ _2249_ _2245_ _2246_ VSS VSS VCC VCC _2250_ sky130_fd_sc_hd__o32a_1
X_3648_ net443 _1527_ _1530_ net733 VSS VSS VCC VCC _1531_ sky130_fd_sc_hd__a211o_1
X_3579_ u_bits.i_op2\[11\] net695 net350 _1465_ VSS VSS VCC VCC _1466_ sky130_fd_sc_hd__o211a_1
X_5318_ clknet_leaf_89_i_clk _0346_ VSS VSS VCC VCC u_muldiv.divisor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_5249_ clknet_leaf_2_i_clk _0277_ VSS VSS VCC VCC u_muldiv.o_div\[26\] sky130_fd_sc_hd__dfxtp_1
X_2950_ net729 _0918_ _0919_ net575 VSS VSS VCC VCC net261 sky130_fd_sc_hd__a211oi_4
X_2881_ net686 net689 net692 net694 net644 net634 VSS VSS VCC VCC _0853_ sky130_fd_sc_hd__mux4_1
X_4620_ u_muldiv.dividend\[7\] net325 net376 _2179_ VSS VSS VCC VCC _0320_
+ sky130_fd_sc_hd__a31o_1
X_4551_ net474 _2115_ _2116_ net438 VSS VSS VCC VCC _2117_ sky130_fd_sc_hd__o31a_1
X_3502_ net456 _1319_ VSS VSS VCC VCC _1394_ sky130_fd_sc_hd__or2_1
X_4482_ _2081_ u_muldiv.quotient_msk\[25\] net433 VSS VSS VCC VCC _2086_ sky130_fd_sc_hd__mux2_1
X_3433_ net412 _1324_ _1326_ _1328_ VSS VSS VCC VCC _1329_ sky130_fd_sc_hd__or4_1
X_3364_ net573 _1213_ _1214_ net565 VSS VSS VCC VCC net311 sky130_fd_sc_hd__a211o_4
X_5103_ clknet_leaf_177_i_clk _0136_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[18\]
+ sky130_fd_sc_hd__dfxtp_2
X_3295_ _0928_ _0970_ _1208_ VSS VSS VCC VCC _1225_ sky130_fd_sc_hd__and3_1
X_5034_ clknet_leaf_22_i_clk _0067_ VSS VSS VCC VCC u_bits.i_op2\[23\] sky130_fd_sc_hd__dfxtp_2
X_4818_ net662 _2358_ VSS VSS VCC VCC _2360_ sky130_fd_sc_hd__nor2_1
X_4749_ u_muldiv.dividend\[18\] net462 _2262_ u_muldiv.dividend\[19\] vssd1 vssd1
+ vccd1 vccd1 _2297_ sky130_fd_sc_hd__o31a_1
Xinput103 i_op2[4] VSS VSS VCC VCC net103 sky130_fd_sc_hd__buf_6
Xinput114 i_pc_next[15] VSS VSS VCC VCC net114 sky130_fd_sc_hd__clkbuf_1
Xinput125 i_pc_target[11] VSS VSS VCC VCC net125 sky130_fd_sc_hd__clkbuf_1
Xinput136 i_pc_target[7] VSS VSS VCC VCC net136 sky130_fd_sc_hd__buf_4
Xinput147 i_reg_data2[12] VSS VSS VCC VCC net147 sky130_fd_sc_hd__clkbuf_1
Xinput158 i_reg_data2[22] VSS VSS VCC VCC net158 sky130_fd_sc_hd__clkbuf_1
Xinput169 i_reg_data2[3] VSS VSS VCC VCC net169 sky130_fd_sc_hd__clkbuf_1
X_3080_ net601 _1040_ net327 VSS VSS VCC VCC _1042_ sky130_fd_sc_hd__o21a_1
X_3982_ u_wr_mux.i_reg_data2\[26\] net162 net398 VSS VSS VCC VCC _0144_ sky130_fd_sc_hd__mux2_1
X_2933_ _0801_ _0809_ _0800_ _0803_ net454 net630 VSS VSS VCC VCC _0903_ sky130_fd_sc_hd__mux4_2
X_2864_ net659 net657 net655 net652 net641 net636 VSS VSS VCC VCC _0836_ sky130_fd_sc_hd__mux4_1
X_4603_ net712 net711 net709 _2131_ net374 VSS VSS VCC VCC _2164_ sky130_fd_sc_hd__o41a_1
X_2795_ net601 _0768_ _0766_ VSS VSS VCC VCC _0769_ sky130_fd_sc_hd__a21oi_2
X_4534_ u_muldiv.quotient_msk\[22\] net480 net334 u_muldiv.quotient_msk\[23\] vssd1
+ vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__a22o_1
X_4465_ net319 _2070_ _2072_ VSS VSS VCC VCC _0272_ sky130_fd_sc_hd__a21oi_1
X_3416_ net557 u_muldiv.mul\[1\] net415 net529 _1312_ VSS VSS VCC VCC _1313_
+ sky130_fd_sc_hd__o311a_2
X_4396_ net320 _2017_ u_muldiv.o_div\[7\] VSS VSS VCC VCC _2018_ sky130_fd_sc_hd__a21o_1
X_3347_ net308 u_wr_mux.i_reg_data2\[23\] net562 VSS VSS VCC VCC net294 sky130_fd_sc_hd__mux2_4
X_3278_ _0576_ _1211_ VSS VSS VCC VCC net183 sky130_fd_sc_hd__and2_4
X_5017_ clknet_leaf_27_i_clk _0050_ VSS VSS VCC VCC u_bits.i_op2\[6\] sky130_fd_sc_hd__dfxtp_4
X_2580_ _0460_ _0549_ _0548_ net428 VSS VSS VCC VCC _0555_ sky130_fd_sc_hd__o211ai_1
X_4250_ _1876_ _1877_ VSS VSS VCC VCC _1878_ sky130_fd_sc_hd__nand2_1
X_3201_ net732 net30 _1156_ VSS VSS VCC VCC net269 sky130_fd_sc_hd__o21a_2
X_4181_ u_muldiv.mul\[11\] u_muldiv.mul\[10\] net403 VSS VSS VCC VCC _0225_
+ sky130_fd_sc_hd__mux2_1
X_3132_ net410 _1079_ _1085_ _1091_ VSS VSS VCC VCC _1092_ sky130_fd_sc_hd__or4_1
X_3063_ net427 _1025_ VSS VSS VCC VCC _1026_ sky130_fd_sc_hd__xor2_1
X_3965_ u_wr_mux.i_reg_data2\[9\] net175 net393 VSS VSS VCC VCC _0127_ sky130_fd_sc_hd__mux2_1
X_2916_ _0744_ _0881_ _0886_ VSS VSS VCC VCC _0887_ sky130_fd_sc_hd__a21oi_4
X_3896_ net509 _1703_ VSS VSS VCC VCC _1704_ sky130_fd_sc_hd__and2b_1
X_2847_ net574 _0820_ VSS VSS VCC VCC _0821_ sky130_fd_sc_hd__nor2_2
X_2778_ _0751_ _0752_ VSS VSS VCC VCC _0753_ sky130_fd_sc_hd__nand2_1
X_4517_ u_muldiv.quotient_msk\[5\] net492 net342 u_muldiv.quotient_msk\[6\] vssd1
+ vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__a22o_1
X_4448_ u_muldiv.o_div\[16\] u_muldiv.o_div\[17\] u_muldiv.o_div\[18\] _2050_ vssd1
+ vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__nor4_2
Xfanout601 net602 VSS VSS VCC VCC net601 sky130_fd_sc_hd__clkbuf_4
Xfanout612 net615 VSS VSS VCC VCC net612 sky130_fd_sc_hd__clkbuf_4
Xfanout623 u_bits.i_op2\[2\] VSS VSS VCC VCC net623 sky130_fd_sc_hd__buf_6
Xfanout634 net635 VSS VSS VCC VCC net634 sky130_fd_sc_hd__clkbuf_8
X_4379_ net322 _2002_ _2004_ u_muldiv.o_div\[3\] VSS VSS VCC VCC _0254_ sky130_fd_sc_hd__o22a_1
Xfanout645 net649 VSS VSS VCC VCC net645 sky130_fd_sc_hd__buf_6
Xfanout656 net657 VSS VSS VCC VCC net656 sky130_fd_sc_hd__buf_4
Xfanout667 net668 VSS VSS VCC VCC net667 sky130_fd_sc_hd__clkbuf_4
Xfanout678 u_bits.i_op1\[19\] VSS VSS VCC VCC net678 sky130_fd_sc_hd__buf_6
Xfanout689 u_bits.i_op1\[14\] VSS VSS VCC VCC net689 sky130_fd_sc_hd__buf_8
X_3750_ net685 net52 net398 VSS VSS VCC VCC _0019_ sky130_fd_sc_hd__mux2_1
X_2701_ net516 net524 _0672_ _0673_ VSS VSS VCC VCC _0676_ sky130_fd_sc_hd__o211ai_1
X_3681_ _0807_ _0980_ _1560_ VSS VSS VCC VCC _1561_ sky130_fd_sc_hd__o21ba_1
X_2632_ net648 net554 net705 net540 net425 VSS VSS VCC VCC _0607_ sky130_fd_sc_hd__o2111ai_4
X_5351_ clknet_leaf_87_i_clk _0378_ VSS VSS VCC VCC u_muldiv.dividend\[0\]
+ sky130_fd_sc_hd__dfxtp_4
Xoutput204 net204 VSS VSS VCC VCC o_add[29] sky130_fd_sc_hd__buf_2
X_2563_ net538 net714 VSS VSS VCC VCC _0538_ sky130_fd_sc_hd__and2_1
Xoutput215 net571 VSS VSS VCC VCC o_funct3[0] sky130_fd_sc_hd__buf_2
Xoutput226 net226 VSS VSS VCC VCC o_pc_target[1] sky130_fd_sc_hd__buf_2
Xoutput237 net237 VSS VSS VCC VCC o_rd[2] sky130_fd_sc_hd__buf_2
Xoutput248 net248 VSS VSS VCC VCC o_result[12] sky130_fd_sc_hd__buf_2
X_4302_ u_muldiv.divisor\[23\] u_muldiv.dividend\[23\] VSS VSS VCC VCC _1930_
+ sky130_fd_sc_hd__nand2b_1
Xoutput259 net259 VSS VSS VCC VCC o_result[22] sky130_fd_sc_hd__buf_2
X_5282_ clknet_leaf_2_i_clk _0310_ VSS VSS VCC VCC u_muldiv.quotient_msk\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_2494_ net671 u_muldiv.add_prev\[22\] net531 VSS VSS VCC VCC _0469_ sky130_fd_sc_hd__mux2_1
X_4233_ u_muldiv.divisor\[2\] _0442_ _1858_ _1860_ VSS VSS VCC VCC _1861_
+ sky130_fd_sc_hd__o211ai_2
X_4164_ net550 net499 net200 VSS VSS VCC VCC _0208_ sky130_fd_sc_hd__o21a_1
X_3115_ u_muldiv.o_div\[29\] net365 _0760_ u_muldiv.mul\[29\] _1074_ vssd1 vssd1 vccd1
+ vccd1 _1075_ sky130_fd_sc_hd__a221o_1
X_4095_ u_muldiv.divisor\[52\] net484 net335 u_muldiv.divisor\[53\] _1802_ vssd1 vssd1
+ vccd1 vccd1 _0172_ sky130_fd_sc_hd__a221o_1
X_3046_ _0852_ net624 net452 _1008_ VSS VSS VCC VCC _1010_ sky130_fd_sc_hd__o211a_1
X_4997_ clknet_leaf_48_i_clk _0030_ VSS VSS VCC VCC u_bits.i_op1\[27\] sky130_fd_sc_hd__dfxtp_4
X_3948_ net559 net42 net395 VSS VSS VCC VCC _0111_ sky130_fd_sc_hd__mux2_1
X_3879_ net584 net586 net546 VSS VSS VCC VCC _1691_ sky130_fd_sc_hd__mux2_1
Xfanout420 net422 VSS VSS VCC VCC net420 sky130_fd_sc_hd__buf_6
Xfanout431 _0457_ VSS VSS VCC VCC net431 sky130_fd_sc_hd__buf_6
Xfanout442 net444 VSS VSS VCC VCC net442 sky130_fd_sc_hd__buf_6
Xfanout453 net455 VSS VSS VCC VCC net453 sky130_fd_sc_hd__buf_4
Xfanout464 u_muldiv.dividend\[1\] VSS VSS VCC VCC net464 sky130_fd_sc_hd__buf_4
Xfanout475 net476 VSS VSS VCC VCC net475 sky130_fd_sc_hd__clkbuf_4
Xfanout486 net487 VSS VSS VCC VCC net486 sky130_fd_sc_hd__buf_2
Xfanout497 net498 VSS VSS VCC VCC net497 sky130_fd_sc_hd__clkbuf_4
X_4920_ u_muldiv.divisor\[27\] net475 net332 u_muldiv.divisor\[28\] vssd1 vssd1 vccd1
+ vccd1 _0372_ sky130_fd_sc_hd__a22o_1
X_4851_ _2388_ net370 net656 net466 VSS VSS VCC VCC _2390_ sky130_fd_sc_hd__a31o_1
X_3802_ net602 net725 _1633_ _1632_ VSS VSS VCC VCC _0048_ sky130_fd_sc_hd__o22a_1
X_4782_ _1928_ _2326_ net467 VSS VSS VCC VCC _2327_ sky130_fd_sc_hd__o21ai_1
X_3733_ net39 net180 VSS VSS VCC VCC _1609_ sky130_fd_sc_hd__nand2b_1
X_3664_ net462 net420 net368 u_muldiv.o_div\[17\] VSS VSS VCC VCC _1545_ sky130_fd_sc_hd__a22oi_4
X_2615_ net710 u_muldiv.add_prev\[4\] net539 VSS VSS VCC VCC _0590_ sky130_fd_sc_hd__mux2_1
X_3595_ net593 net694 VSS VSS VCC VCC _1481_ sky130_fd_sc_hd__nand2_1
X_2546_ net535 _0428_ _0520_ VSS VSS VCC VCC _0521_ sky130_fd_sc_hd__o21ai_1
X_5334_ clknet_leaf_147_i_clk _0362_ VSS VSS VCC VCC u_muldiv.divisor\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_130_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_130_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5265_ clknet_leaf_120_i_clk _0293_ VSS VSS VCC VCC u_muldiv.quotient_msk\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2477_ u_muldiv.o_div\[8\] VSS VSS VCC VCC _0452_ sky130_fd_sc_hd__inv_2
X_4216_ u_muldiv.dividend\[9\] u_muldiv.divisor\[9\] VSS VSS VCC VCC _1844_
+ sky130_fd_sc_hd__nand2b_1
X_5196_ clknet_4_9__leaf_i_clk _0228_ VSS VSS VCC VCC u_muldiv.mul\[13\] sky130_fd_sc_hd__dfxtp_1
X_4147_ net555 net500 net213 VSS VSS VCC VCC _0191_ sky130_fd_sc_hd__o21a_1
X_4078_ _1787_ net380 net588 net329 VSS VSS VCC VCC _1789_ sky130_fd_sc_hd__a31o_1
X_3029_ net516 net523 _0992_ VSS VSS VCC VCC _0994_ sky130_fd_sc_hd__o21ai_1
X_3380_ _1277_ _1272_ net607 VSS VSS VCC VCC _1278_ sky130_fd_sc_hd__mux2_1
X_5050_ clknet_leaf_81_i_clk _0083_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_4001_ net640 net626 net378 VSS VSS VCC VCC _1728_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_77_i_clk clknet_4_13__leaf_i_clk VSS VSS VCC VCC clknet_leaf_77_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4903_ u_muldiv.divisor\[10\] net490 net338 u_muldiv.divisor\[11\] vssd1 vssd1 vccd1
+ vccd1 _0355_ sky130_fd_sc_hd__a22o_1
X_4834_ _2371_ _2374_ _2373_ net433 VSS VSS VCC VCC _2375_ sky130_fd_sc_hd__a22o_1
X_4765_ net481 _2311_ _2306_ net317 VSS VSS VCC VCC _2312_ sky130_fd_sc_hd__o211a_1
X_3716_ net730 _1593_ net576 VSS VSS VCC VCC _1594_ sky130_fd_sc_hd__a21oi_1
X_4696_ net693 net690 _2227_ net372 net688 VSS VSS VCC VCC _2249_ sky130_fd_sc_hd__o311a_1
X_3647_ net556 u_muldiv.mul\[15\] net415 net528 _1529_ VSS VSS VCC VCC _1530_
+ sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_15_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_15_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3578_ net566 _0438_ net594 VSS VSS VCC VCC _1465_ sky130_fd_sc_hd__or3b_1
X_5317_ clknet_leaf_89_i_clk _0345_ VSS VSS VCC VCC u_muldiv.divisor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2529_ _0502_ _0503_ VSS VSS VCC VCC _0504_ sky130_fd_sc_hd__nand2_1
X_5248_ clknet_leaf_3_i_clk _0276_ VSS VSS VCC VCC u_muldiv.o_div\[25\] sky130_fd_sc_hd__dfxtp_2
X_5179_ clknet_4_7__leaf_i_clk _0211_ VSS VSS VCC VCC u_muldiv.add_prev\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_2880_ net696 net698 net700 net703 net644 net635 VSS VSS VCC VCC _0852_ sky130_fd_sc_hd__mux4_2
X_4550_ net461 net374 net717 VSS VSS VCC VCC _2116_ sky130_fd_sc_hd__a21oi_1
X_3501_ _1393_ u_pc_sel.i_pc_next\[5\] net575 VSS VSS VCC VCC net272 sky130_fd_sc_hd__mux2_1
X_4481_ _2081_ net475 u_muldiv.o_div\[25\] net383 VSS VSS VCC VCC _2085_ sky130_fd_sc_hd__a31o_1
X_3432_ net621 net715 net350 _1327_ VSS VSS VCC VCC _1328_ sky130_fd_sc_hd__o211a_1
Xclkbuf_4_5__f_i_clk clknet_2_1_0_i_clk VSS VSS VCC VCC clknet_4_5__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3363_ u_wr_mux.i_reg_data2\[15\] _0764_ _1265_ VSS VSS VCC VCC net303 sky130_fd_sc_hd__a21o_4
X_5102_ clknet_leaf_34_i_clk _0135_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_3294_ _1223_ _1140_ VSS VSS VCC VCC _1224_ sky130_fd_sc_hd__nand2_1
X_5033_ clknet_leaf_28_i_clk _0066_ VSS VSS VCC VCC u_bits.i_op2\[22\] sky130_fd_sc_hd__dfxtp_4
X_4817_ net667 net664 _2338_ net369 net662 VSS VSS VCC VCC _2359_ sky130_fd_sc_hd__o311a_1
X_4748_ _1912_ _2295_ VSS VSS VCC VCC _2296_ sky130_fd_sc_hd__xor2_1
X_4679_ _1894_ _1895_ _2225_ net470 VSS VSS VCC VCC _2233_ sky130_fd_sc_hd__o31a_1
Xinput104 i_op2[5] VSS VSS VCC VCC net104 sky130_fd_sc_hd__clkbuf_1
Xinput115 i_pc_next[1] VSS VSS VCC VCC net115 sky130_fd_sc_hd__clkbuf_1
Xinput126 i_pc_target[12] VSS VSS VCC VCC net126 sky130_fd_sc_hd__clkbuf_2
Xinput137 i_pc_target[8] VSS VSS VCC VCC net137 sky130_fd_sc_hd__buf_8
Xinput148 i_reg_data2[13] VSS VSS VCC VCC net148 sky130_fd_sc_hd__clkbuf_1
Xinput159 i_reg_data2[23] VSS VSS VCC VCC net159 sky130_fd_sc_hd__dlymetal6s2s_1
X_3981_ u_wr_mux.i_reg_data2\[25\] net161 net396 VSS VSS VCC VCC _0143_ sky130_fd_sc_hd__mux2_1
X_2932_ _0809_ _0803_ net630 VSS VSS VCC VCC _0902_ sky130_fd_sc_hd__mux2_1
X_2863_ net654 net652 net638 VSS VSS VCC VCC _0835_ sky130_fd_sc_hd__mux2_1
X_4602_ _1865_ _1849_ _1850_ _1867_ _1847_ VSS VSS VCC VCC _2163_ sky130_fd_sc_hd__a311o_1
X_2794_ net650 u_bits.i_sra VSS VSS VCC VCC _0768_ sky130_fd_sc_hd__nand2_1
X_4533_ u_muldiv.quotient_msk\[21\] net488 net341 u_muldiv.quotient_msk\[22\] vssd1
+ vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__a22o_1
X_4464_ net319 _2071_ u_muldiv.o_div\[21\] VSS VSS VCC VCC _2072_ sky130_fd_sc_hd__a21oi_1
X_3415_ u_muldiv.o_div\[1\] net367 net359 _1311_ VSS VSS VCC VCC _1312_ sky130_fd_sc_hd__a211o_1
X_4395_ u_muldiv.quotient_msk\[7\] net438 _2013_ VSS VSS VCC VCC _2017_ sky130_fd_sc_hd__a21o_1
X_3346_ net307 u_wr_mux.i_reg_data2\[22\] net563 VSS VSS VCC VCC net293 sky130_fd_sc_hd__mux2_8
X_3277_ _0574_ _0575_ _0573_ VSS VSS VCC VCC _1211_ sky130_fd_sc_hd__or3_2
X_5016_ clknet_leaf_34_i_clk _0049_ VSS VSS VCC VCC u_bits.i_op2\[5\] sky130_fd_sc_hd__dfxtp_4
X_3200_ net575 _1155_ VSS VSS VCC VCC _1156_ sky130_fd_sc_hd__nor2_4
X_4180_ u_muldiv.mul\[10\] u_muldiv.mul\[9\] net403 VSS VSS VCC VCC _0224_
+ sky130_fd_sc_hd__mux2_1
X_3131_ net601 _0814_ _1082_ _1090_ VSS VSS VCC VCC _1091_ sky130_fd_sc_hd__a31o_1
X_3062_ net445 u_bits.i_op2\[28\] _0464_ net657 VSS VSS VCC VCC _1025_ sky130_fd_sc_hd__a22o_1
X_3964_ u_wr_mux.i_reg_data2\[8\] net174 net396 VSS VSS VCC VCC _0126_ sky130_fd_sc_hd__mux2_1
X_2915_ _0528_ _0879_ _0884_ _0883_ VSS VSS VCC VCC _0886_ sky130_fd_sc_hd__a211o_1
X_3895_ u_bits.i_op2\[29\] u_bits.i_op2\[27\] net550 VSS VSS VCC VCC _1703_
+ sky130_fd_sc_hd__mux2_1
X_2846_ _0761_ _0819_ net735 VSS VSS VCC VCC _0820_ sky130_fd_sc_hd__a21oi_1
X_2777_ _0750_ _0473_ VSS VSS VCC VCC _0752_ sky130_fd_sc_hd__nand2_1
X_4516_ u_muldiv.quotient_msk\[4\] net496 net342 u_muldiv.quotient_msk\[5\] vssd1
+ vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__a22o_1
X_4447_ u_muldiv.o_div\[16\] u_muldiv.o_div\[17\] _2050_ VSS VSS VCC VCC _2058_
+ sky130_fd_sc_hd__or3_2
Xfanout602 net603 VSS VSS VCC VCC net602 sky130_fd_sc_hd__clkbuf_4
Xfanout613 net614 VSS VSS VCC VCC net613 sky130_fd_sc_hd__buf_2
Xfanout624 u_bits.i_op2\[2\] VSS VSS VCC VCC net624 sky130_fd_sc_hd__buf_8
Xfanout635 net636 VSS VSS VCC VCC net635 sky130_fd_sc_hd__buf_2
X_4378_ net325 net376 _2003_ VSS VSS VCC VCC _2004_ sky130_fd_sc_hd__a21oi_1
Xfanout646 net647 VSS VSS VCC VCC net646 sky130_fd_sc_hd__buf_6
Xfanout657 u_bits.i_op1\[28\] VSS VSS VCC VCC net657 sky130_fd_sc_hd__clkbuf_8
X_3329_ net549 net499 VSS VSS VCC VCC _1256_ sky130_fd_sc_hd__or2_4
Xfanout668 net669 VSS VSS VCC VCC net668 sky130_fd_sc_hd__buf_2
Xfanout679 net680 VSS VSS VCC VCC net679 sky130_fd_sc_hd__clkbuf_4
X_2700_ net516 net523 _0672_ _0673_ VSS VSS VCC VCC _0675_ sky130_fd_sc_hd__o211a_1
X_3680_ net613 _0978_ _1325_ net607 net409 VSS VSS VCC VCC _1560_ sky130_fd_sc_hd__a221o_1
X_2631_ _0582_ _0583_ _0604_ VSS VSS VCC VCC _0606_ sky130_fd_sc_hd__a21o_1
X_5350_ clknet_leaf_93_i_clk _0377_ VSS VSS VCC VCC u_muldiv.o_div\[0\] sky130_fd_sc_hd__dfxtp_2
Xoutput205 net205 VSS VSS VCC VCC o_add[2] sky130_fd_sc_hd__buf_2
X_2562_ net447 net617 VSS VSS VCC VCC _0537_ sky130_fd_sc_hd__nand2_1
Xoutput216 net563 VSS VSS VCC VCC o_funct3[1] sky130_fd_sc_hd__buf_2
Xoutput227 net227 VSS VSS VCC VCC o_pc_target[2] sky130_fd_sc_hd__buf_2
Xoutput238 net238 VSS VSS VCC VCC o_rd[3] sky130_fd_sc_hd__buf_2
X_4301_ u_muldiv.divisor\[23\] u_muldiv.dividend\[23\] VSS VSS VCC VCC _1929_
+ sky130_fd_sc_hd__and2b_1
Xoutput249 net249 VSS VSS VCC VCC o_result[13] sky130_fd_sc_hd__buf_2
X_5281_ clknet_leaf_178_i_clk _0309_ VSS VSS VCC VCC u_muldiv.quotient_msk\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_2493_ _0465_ _0466_ net427 VSS VSS VCC VCC _0468_ sky130_fd_sc_hd__o21ai_2
X_4232_ u_muldiv.divisor\[0\] _0440_ net464 _0418_ VSS VSS VCC VCC _1860_
+ sky130_fd_sc_hd__o2bb2ai_1
X_4163_ net549 net499 net199 VSS VSS VCC VCC _0207_ sky130_fd_sc_hd__o21a_1
X_3114_ net565 net558 u_muldiv.dividend\[29\] net443 VSS VSS VCC VCC _1074_
+ sky130_fd_sc_hd__a31o_2
X_4094_ u_bits.i_op2\[21\] _1800_ _1801_ VSS VSS VCC VCC _1802_ sky130_fd_sc_hd__o21ba_1
X_3045_ net623 _0852_ _1008_ VSS VSS VCC VCC _1009_ sky130_fd_sc_hd__o21ai_1
X_4996_ clknet_leaf_133_i_clk _0029_ VSS VSS VCC VCC u_bits.i_op1\[26\] sky130_fd_sc_hd__dfxtp_4
X_3947_ net562 net41 net387 VSS VSS VCC VCC _0110_ sky130_fd_sc_hd__mux2_1
X_3878_ net586 net725 _1690_ _1689_ VSS VSS VCC VCC _0067_ sky130_fd_sc_hd__o22a_1
X_2829_ net458 net688 _0802_ VSS VSS VCC VCC _0803_ sky130_fd_sc_hd__a21oi_1
Xfanout410 net412 VSS VSS VCC VCC net410 sky130_fd_sc_hd__buf_4
Xfanout421 net422 VSS VSS VCC VCC net421 sky130_fd_sc_hd__clkbuf_4
Xfanout432 _0457_ VSS VSS VCC VCC net432 sky130_fd_sc_hd__buf_6
Xfanout443 net444 VSS VSS VCC VCC net443 sky130_fd_sc_hd__buf_4
Xfanout454 net455 VSS VSS VCC VCC net454 sky130_fd_sc_hd__buf_4
Xfanout465 net466 VSS VSS VCC VCC net465 sky130_fd_sc_hd__buf_6
Xfanout476 net487 VSS VSS VCC VCC net476 sky130_fd_sc_hd__buf_4
Xfanout487 u_muldiv.i_on_end VSS VSS VCC VCC net487 sky130_fd_sc_hd__buf_6
Xfanout498 u_muldiv.i_on_end VSS VSS VCC VCC net498 sky130_fd_sc_hd__buf_2
X_4850_ _2388_ net370 net656 VSS VSS VCC VCC _2389_ sky130_fd_sc_hd__a21oi_1
X_3801_ net505 net103 net719 VSS VSS VCC VCC _1633_ sky130_fd_sc_hd__a21o_1
X_4781_ _1940_ _1925_ _1942_ VSS VSS VCC VCC _2326_ sky130_fd_sc_hd__o21bai_1
X_3732_ net39 net180 VSS VSS VCC VCC _1608_ sky130_fd_sc_hd__and2b_4
X_3663_ net729 net13 _1544_ VSS VSS VCC VCC net252 sky130_fd_sc_hd__o21a_1
X_2614_ net429 _0585_ _0586_ VSS VSS VCC VCC _0589_ sky130_fd_sc_hd__and3_1
X_3594_ _1041_ net604 _0766_ _1479_ VSS VSS VCC VCC _1480_ sky130_fd_sc_hd__a211oi_1
X_5333_ clknet_leaf_144_i_clk _0361_ VSS VSS VCC VCC u_muldiv.divisor\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_2545_ net647 net552 net685 net535 net424 VSS VSS VCC VCC _0520_ sky130_fd_sc_hd__o2111ai_4
X_5264_ clknet_leaf_119_i_clk _0292_ VSS VSS VCC VCC u_muldiv.quotient_msk\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2476_ net491 VSS VSS VCC VCC _0451_ sky130_fd_sc_hd__inv_2
X_4215_ u_muldiv.divisor\[30\] _0447_ VSS VSS VCC VCC _1843_ sky130_fd_sc_hd__nor2_1
X_5195_ clknet_leaf_111_i_clk _0227_ VSS VSS VCC VCC u_muldiv.mul\[12\] sky130_fd_sc_hd__dfxtp_1
X_4146_ _1173_ _1174_ net401 VSS VSS VCC VCC _0190_ sky130_fd_sc_hd__and3_1
X_4077_ _1787_ net380 net588 VSS VSS VCC VCC _1788_ sky130_fd_sc_hd__a21oi_1
X_3028_ net533 net659 _0463_ _0991_ net427 VSS VSS VCC VCC _0993_ sky130_fd_sc_hd__a311o_1
X_4979_ clknet_leaf_51_i_clk _0012_ VSS VSS VCC VCC u_bits.i_op1\[9\] sky130_fd_sc_hd__dfxtp_1
X_4000_ u_muldiv.divisor\[32\] net478 net333 u_muldiv.divisor\[33\] _1727_ vssd1 vssd1
+ vccd1 vccd1 _0152_ sky130_fd_sc_hd__a221o_1
X_4902_ u_muldiv.divisor\[9\] net494 net339 u_muldiv.divisor\[10\] vssd1 vssd1 vccd1
+ vccd1 _0354_ sky130_fd_sc_hd__a22o_1
X_4833_ u_muldiv.dividend\[26\] u_muldiv.dividend\[25\] _2345_ net476 vssd1 vssd1
+ vccd1 vccd1 _2374_ sky130_fd_sc_hd__o31a_1
X_4764_ net467 _2310_ _2308_ VSS VSS VCC VCC _2311_ sky130_fd_sc_hd__o21ai_1
X_3715_ net444 _1582_ _1583_ _1592_ VSS VSS VCC VCC _1593_ sky130_fd_sc_hd__o31ai_1
X_4695_ net688 _2247_ VSS VSS VCC VCC _2248_ sky130_fd_sc_hd__nor2_1
X_3646_ u_muldiv.dividend\[15\] net421 net358 _1528_ VSS VSS VCC VCC _1529_
+ sky130_fd_sc_hd__a211o_1
X_3577_ net578 u_pc_sel.i_pc_next\[10\] _1463_ _1464_ VSS VSS VCC VCC net246
+ sky130_fd_sc_hd__a22o_4
X_5316_ clknet_leaf_17_i_clk _0344_ VSS VSS VCC VCC u_muldiv.dividend\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_2528_ _0500_ _0501_ net427 VSS VSS VCC VCC _0503_ sky130_fd_sc_hd__a21o_1
X_5247_ clknet_4_3__leaf_i_clk _0275_ VSS VSS VCC VCC u_muldiv.o_div\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_2459_ net559 VSS VSS VCC VCC _0434_ sky130_fd_sc_hd__inv_4
X_5178_ clknet_4_7__leaf_i_clk _0210_ VSS VSS VCC VCC u_muldiv.add_prev\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_4129_ _1827_ net378 net581 net329 VSS VSS VCC VCC _1829_ sky130_fd_sc_hd__a31o_1
X_3500_ _1392_ net33 net735 VSS VSS VCC VCC _1393_ sky130_fd_sc_hd__mux2_2
X_4480_ u_muldiv.o_div\[24\] _2084_ net317 VSS VSS VCC VCC _0275_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_144_i_clk clknet_4_8__leaf_i_clk VSS VSS VCC VCC clknet_leaf_144_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3431_ net457 net565 net715 VSS VSS VCC VCC _1327_ sky130_fd_sc_hd__or3b_1
X_3362_ net216 u_wr_mux.i_reg_data2\[31\] net417 net308 VSS VSS VCC VCC _1265_
+ sky130_fd_sc_hd__a22o_1
X_5101_ clknet_leaf_135_i_clk _0134_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_3293_ _1109_ _1110_ _1002_ _1073_ VSS VSS VCC VCC _1223_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_159_i_clk clknet_4_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_159_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5032_ clknet_leaf_27_i_clk _0065_ VSS VSS VCC VCC u_bits.i_op2\[21\] sky130_fd_sc_hd__dfxtp_4
X_4816_ net667 net664 _2338_ net369 VSS VSS VCC VCC _2358_ sky130_fd_sc_hd__o31a_1
X_4747_ u_muldiv.divisor\[18\] _0450_ _2286_ VSS VSS VCC VCC _2295_ sky130_fd_sc_hd__o21ai_1
X_4678_ _1895_ _2225_ _1894_ VSS VSS VCC VCC _2232_ sky130_fd_sc_hd__o21ai_1
X_3629_ net356 _1204_ _1512_ VSS VSS VCC VCC _1513_ sky130_fd_sc_hd__o21ai_1
Xinput105 i_op2[6] VSS VSS VCC VCC net105 sky130_fd_sc_hd__buf_6
Xinput116 i_pc_next[2] VSS VSS VCC VCC net116 sky130_fd_sc_hd__buf_2
Xinput127 i_pc_target[13] VSS VSS VCC VCC net127 sky130_fd_sc_hd__buf_8
Xinput138 i_pc_target[9] VSS VSS VCC VCC net138 sky130_fd_sc_hd__clkbuf_4
Xinput149 i_reg_data2[14] VSS VSS VCC VCC net149 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_61_i_clk clknet_4_7__leaf_i_clk VSS VSS VCC VCC clknet_leaf_61_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_76_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_76_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_14_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_14_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3980_ u_wr_mux.i_reg_data2\[24\] net160 net389 VSS VSS VCC VCC _0142_ sky130_fd_sc_hd__mux2_1
X_2931_ net603 _0814_ VSS VSS VCC VCC _0901_ sky130_fd_sc_hd__nand2_2
X_2862_ u_muldiv.mul\[55\] net363 net357 u_muldiv.mul\[23\] _0833_ vssd1 vssd1 vccd1
+ vccd1 _0834_ sky130_fd_sc_hd__a221o_2
X_4601_ _2160_ _2161_ net438 VSS VSS VCC VCC _2162_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_29_i_clk clknet_4_4__leaf_i_clk VSS VSS VCC VCC clknet_leaf_29_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2793_ net650 u_bits.i_sra VSS VSS VCC VCC _0767_ sky130_fd_sc_hd__and2_1
X_4532_ u_muldiv.quotient_msk\[20\] net489 net341 u_muldiv.quotient_msk\[21\] vssd1
+ vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__a22o_1
X_4463_ _2066_ u_muldiv.quotient_msk\[21\] net437 VSS VSS VCC VCC _2071_ sky130_fd_sc_hd__mux2_1
X_3414_ net568 net557 net464 u_muldiv.mul\[33\] net361 VSS VSS VCC VCC _1311_
+ sky130_fd_sc_hd__a32o_1
X_4394_ u_muldiv.o_div\[7\] _2013_ net473 net493 VSS VSS VCC VCC _2016_ sky130_fd_sc_hd__o2bb2a_1
X_3345_ net306 u_wr_mux.i_reg_data2\[21\] net565 VSS VSS VCC VCC net292 sky130_fd_sc_hd__mux2_4
X_3276_ _0745_ _0748_ VSS VSS VCC VCC net195 sky130_fd_sc_hd__xor2_4
X_5015_ clknet_leaf_15_i_clk _0048_ VSS VSS VCC VCC u_bits.i_op2\[4\] sky130_fd_sc_hd__dfxtp_4
X_3130_ _1087_ net611 _1089_ VSS VSS VCC VCC _1090_ sky130_fd_sc_hd__a21oi_1
X_3061_ net732 net25 _1024_ VSS VSS VCC VCC net264 sky130_fd_sc_hd__o21a_1
X_3963_ net308 net173 net390 VSS VSS VCC VCC _0125_ sky130_fd_sc_hd__mux2_1
X_2914_ _0528_ _0879_ _0884_ _0883_ VSS VSS VCC VCC _0885_ sky130_fd_sc_hd__a211oi_2
X_3894_ net582 net723 _1702_ _1701_ VSS VSS VCC VCC _0071_ sky130_fd_sc_hd__o22a_1
X_2845_ _0422_ _0818_ net197 net355 net527 VSS VSS VCC VCC _0819_ sky130_fd_sc_hd__a221o_1
X_2776_ _0749_ _0745_ _0489_ _0474_ VSS VSS VCC VCC _0751_ sky130_fd_sc_hd__o211ai_1
X_4515_ u_muldiv.quotient_msk\[3\] net496 net342 u_muldiv.quotient_msk\[4\] vssd1
+ vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__a22o_1
X_4446_ net322 _2055_ _2057_ u_muldiv.o_div\[17\] VSS VSS VCC VCC _0268_ sky130_fd_sc_hd__o22a_1
Xfanout603 u_bits.i_op2\[4\] VSS VSS VCC VCC net603 sky130_fd_sc_hd__buf_4
X_4377_ u_muldiv.quotient_msk\[3\] net438 _1999_ VSS VSS VCC VCC _2003_ sky130_fd_sc_hd__a21oi_1
Xfanout614 net615 VSS VSS VCC VCC net614 sky130_fd_sc_hd__buf_4
Xfanout625 net633 VSS VSS VCC VCC net625 sky130_fd_sc_hd__buf_4
Xfanout636 u_bits.i_op2\[1\] VSS VSS VCC VCC net636 sky130_fd_sc_hd__buf_4
Xfanout647 net648 VSS VSS VCC VCC net647 sky130_fd_sc_hd__buf_6
X_3328_ net550 net500 VSS VSS VCC VCC _1255_ sky130_fd_sc_hd__nor2_2
Xfanout658 u_bits.i_op1\[27\] VSS VSS VCC VCC net658 sky130_fd_sc_hd__buf_4
Xfanout669 u_bits.i_op1\[23\] VSS VSS VCC VCC net669 sky130_fd_sc_hd__buf_4
X_3259_ _0736_ _1191_ _0650_ _0661_ VSS VSS VCC VCC _1199_ sky130_fd_sc_hd__o211ai_2
X_2630_ _0582_ _0583_ _0604_ VSS VSS VCC VCC _0605_ sky130_fd_sc_hd__a21oi_2
X_2561_ net448 net714 _0534_ VSS VSS VCC VCC _0536_ sky130_fd_sc_hd__a21oi_1
Xoutput206 net206 VSS VSS VCC VCC o_add[30] sky130_fd_sc_hd__buf_2
Xoutput217 net559 VSS VSS VCC VCC o_funct3[2] sky130_fd_sc_hd__buf_2
X_4300_ _1926_ _1927_ VSS VSS VCC VCC _1928_ sky130_fd_sc_hd__nor2_1
Xoutput228 net228 VSS VSS VCC VCC o_pc_target[3] sky130_fd_sc_hd__buf_2
Xoutput239 net239 VSS VSS VCC VCC o_rd[4] sky130_fd_sc_hd__buf_2
X_5280_ clknet_leaf_178_i_clk _0308_ VSS VSS VCC VCC u_muldiv.quotient_msk\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_2492_ net671 net531 _0463_ _0466_ net430 VSS VSS VCC VCC _0467_ sky130_fd_sc_hd__a311o_1
X_4231_ _0440_ u_muldiv.divisor\[0\] VSS VSS VCC VCC _1859_ sky130_fd_sc_hd__nand2_1
X_4162_ net549 net499 net198 VSS VSS VCC VCC _0206_ sky130_fd_sc_hd__o21a_1
X_3113_ _1073_ VSS VSS VCC VCC net204 sky130_fd_sc_hd__clkinv_4
X_4093_ u_bits.i_op2\[21\] _1800_ net484 net468 VSS VSS VCC VCC _1801_ sky130_fd_sc_hd__a211o_1
X_3044_ net457 _0845_ VSS VSS VCC VCC _1008_ sky130_fd_sc_hd__or2_1
X_4995_ clknet_leaf_164_i_clk _0028_ VSS VSS VCC VCC u_bits.i_op1\[25\] sky130_fd_sc_hd__dfxtp_1
X_3946_ net570 net40 net387 VSS VSS VCC VCC _0109_ sky130_fd_sc_hd__mux2_1
X_3877_ net507 net92 net719 VSS VSS VCC VCC _1690_ sky130_fd_sc_hd__a21o_1
X_2828_ net643 net691 VSS VSS VCC VCC _0802_ sky130_fd_sc_hd__and2_1
X_2759_ _0724_ _0712_ _0725_ VSS VSS VCC VCC _0734_ sky130_fd_sc_hd__a21boi_2
X_4429_ u_muldiv.o_div\[13\] _2035_ u_muldiv.o_div\[14\] VSS VSS VCC VCC _2044_
+ sky130_fd_sc_hd__o21a_1
Xfanout400 _1256_ VSS VSS VCC VCC net400 sky130_fd_sc_hd__buf_8
Xfanout411 net412 VSS VSS VCC VCC net411 sky130_fd_sc_hd__clkbuf_4
Xfanout422 _0754_ VSS VSS VCC VCC net422 sky130_fd_sc_hd__buf_4
Xfanout433 net434 VSS VSS VCC VCC net433 sky130_fd_sc_hd__buf_6
Xfanout444 _0423_ VSS VSS VCC VCC net444 sky130_fd_sc_hd__clkbuf_8
Xfanout455 _0420_ VSS VSS VCC VCC net455 sky130_fd_sc_hd__clkbuf_4
Xfanout466 net467 VSS VSS VCC VCC net466 sky130_fd_sc_hd__clkbuf_8
Xfanout477 net478 VSS VSS VCC VCC net477 sky130_fd_sc_hd__clkbuf_4
Xfanout488 net495 VSS VSS VCC VCC net488 sky130_fd_sc_hd__buf_4
Xfanout499 net500 VSS VSS VCC VCC net499 sky130_fd_sc_hd__buf_6
X_3800_ net505 _1631_ VSS VSS VCC VCC _1632_ sky130_fd_sc_hd__and2b_1
X_4780_ u_muldiv.dividend\[22\] _2280_ _2321_ _0450_ VSS VSS VCC VCC _2325_
+ sky130_fd_sc_hd__and4b_1
X_3731_ net731 net19 _1607_ VSS VSS VCC VCC net258 sky130_fd_sc_hd__o21a_2
X_3662_ net729 _1543_ net576 VSS VSS VCC VCC _1544_ sky130_fd_sc_hd__a21oi_1
X_2613_ _0459_ net425 net539 net711 net431 VSS VSS VCC VCC _0588_ sky130_fd_sc_hd__a41oi_1
X_3593_ _0806_ _1359_ _1363_ _0856_ VSS VSS VCC VCC _1479_ sky130_fd_sc_hd__a22o_1
X_5332_ clknet_leaf_143_i_clk _0360_ VSS VSS VCC VCC u_muldiv.divisor\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_2544_ _0513_ _0514_ _0517_ VSS VSS VCC VCC _0519_ sky130_fd_sc_hd__nand3b_1
X_5263_ clknet_leaf_119_i_clk _0291_ VSS VSS VCC VCC u_muldiv.quotient_msk\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_2475_ u_muldiv.dividend\[18\] VSS VSS VCC VCC _0450_ sky130_fd_sc_hd__inv_2
X_4214_ op_cnt\[5\] _1841_ _1842_ VSS VSS VCC VCC _0251_ sky130_fd_sc_hd__o21ba_1
X_5194_ clknet_leaf_111_i_clk _0226_ VSS VSS VCC VCC u_muldiv.mul\[11\] sky130_fd_sc_hd__dfxtp_1
X_4145_ _1172_ _1176_ net401 VSS VSS VCC VCC _0189_ sky130_fd_sc_hd__and3_1
X_4076_ net591 net590 net589 _1775_ VSS VSS VCC VCC _1787_ sky130_fd_sc_hd__or4_2
X_3027_ net533 net659 _0463_ _0991_ VSS VSS VCC VCC _0992_ sky130_fd_sc_hd__a31o_1
X_4978_ clknet_leaf_82_i_clk _0011_ VSS VSS VCC VCC u_bits.i_op1\[8\] sky130_fd_sc_hd__dfxtp_1
X_3929_ net179 net513 VSS VSS VCC VCC _1716_ sky130_fd_sc_hd__nand2b_1
X_4901_ u_muldiv.divisor\[8\] net494 net339 u_muldiv.divisor\[9\] vssd1 vssd1 vccd1
+ vccd1 _0353_ sky130_fd_sc_hd__a22o_1
X_4832_ _2367_ net465 _2366_ _2369_ _2370_ VSS VSS VCC VCC _2373_ sky130_fd_sc_hd__a32o_1
X_4763_ net675 _2309_ VSS VSS VCC VCC _2310_ sky130_fd_sc_hd__xnor2_1
X_3714_ net195 net354 net530 _1591_ VSS VSS VCC VCC _1592_ sky130_fd_sc_hd__a211o_1
X_4694_ net693 net690 _2227_ net372 VSS VSS VCC VCC _2247_ sky130_fd_sc_hd__o31a_1
X_3645_ net441 net413 u_muldiv.mul\[47\] u_muldiv.o_div\[15\] net366 vssd1 vssd1 vccd1
+ vccd1 _1528_ sky130_fd_sc_hd__a32o_1
X_3576_ net7 net732 net578 VSS VSS VCC VCC _1464_ sky130_fd_sc_hd__o21ba_1
X_2527_ net516 net523 _0500_ _0501_ VSS VSS VCC VCC _0502_ sky130_fd_sc_hd__o211ai_1
X_5315_ clknet_4_1__leaf_i_clk _0343_ VSS VSS VCC VCC u_muldiv.dividend\[30\]
+ sky130_fd_sc_hd__dfxtp_2
X_2458_ net2 VSS VSS VCC VCC _0433_ sky130_fd_sc_hd__inv_2
X_5246_ clknet_leaf_158_i_clk _0274_ VSS VSS VCC VCC u_muldiv.o_div\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_5177_ clknet_leaf_58_i_clk _0209_ VSS VSS VCC VCC u_muldiv.add_prev\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_4128_ _1827_ net378 net581 VSS VSS VCC VCC _1828_ sky130_fd_sc_hd__a21oi_1
X_4059_ u_muldiv.divisor\[45\] net485 net335 u_muldiv.divisor\[46\] _1773_ vssd1 vssd1
+ vccd1 vccd1 _0165_ sky130_fd_sc_hd__a221o_1
X_3430_ _0910_ _1325_ VSS VSS VCC VCC _1326_ sky130_fd_sc_hd__nor2_1
X_3361_ u_wr_mux.i_reg_data2\[14\] _0764_ _1264_ VSS VSS VCC VCC net302 sky130_fd_sc_hd__a21o_1
X_5100_ clknet_leaf_78_i_clk _0133_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_3292_ net203 _1201_ _0832_ _1210_ VSS VSS VCC VCC _1222_ sky130_fd_sc_hd__nand4b_1
X_5031_ clknet_leaf_30_i_clk _0064_ VSS VSS VCC VCC u_bits.i_op2\[20\] sky130_fd_sc_hd__dfxtp_4
X_4815_ _1947_ _2355_ _2356_ VSS VSS VCC VCC _2357_ sky130_fd_sc_hd__a21oi_1
X_4746_ u_muldiv.dividend\[18\] net326 net377 _2294_ VSS VSS VCC VCC _0331_
+ sky130_fd_sc_hd__a31o_1
X_4677_ u_muldiv.dividend\[12\] net324 net375 _2231_ VSS VSS VCC VCC _0325_
+ sky130_fd_sc_hd__a31o_1
X_3628_ net412 _1508_ _1511_ _1507_ net520 VSS VSS VCC VCC _1512_ sky130_fd_sc_hd__a221o_1
X_3559_ net559 u_muldiv.mul\[9\] net414 net529 VSS VSS VCC VCC _1448_ sky130_fd_sc_hd__o31a_1
Xinput106 i_op2[7] VSS VSS VCC VCC net106 sky130_fd_sc_hd__buf_6
Xinput117 i_pc_next[3] VSS VSS VCC VCC net117 sky130_fd_sc_hd__clkbuf_1
Xinput128 i_pc_target[14] VSS VSS VCC VCC net128 sky130_fd_sc_hd__clkbuf_2
Xinput139 i_rd[0] VSS VSS VCC VCC net139 sky130_fd_sc_hd__clkbuf_2
X_5229_ clknet_leaf_114_i_clk _0257_ VSS VSS VCC VCC u_muldiv.o_div\[6\] sky130_fd_sc_hd__dfxtp_2
X_2930_ net628 _0791_ _0897_ _0899_ net613 VSS VSS VCC VCC _0900_ sky130_fd_sc_hd__o32a_2
X_2861_ u_muldiv.dividend\[23\] net419 net364 u_muldiv.o_div\[23\] net442 vssd1 vssd1
+ vccd1 vccd1 _0833_ sky130_fd_sc_hd__a221o_1
X_4600_ u_muldiv.dividend\[5\] _2136_ _0444_ _0443_ VSS VSS VCC VCC _2161_
+ sky130_fd_sc_hd__nand4b_4
X_2792_ net564 net440 net573 VSS VSS VCC VCC _0766_ sky130_fd_sc_hd__or3b_2
X_4531_ u_muldiv.quotient_msk\[19\] net490 net338 u_muldiv.quotient_msk\[20\] vssd1
+ vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__a22o_1
X_4462_ _2066_ u_muldiv.o_div\[21\] net488 net385 VSS VSS VCC VCC _2070_ sky130_fd_sc_hd__a31o_1
X_3413_ _0422_ net194 _1309_ net443 VSS VSS VCC VCC _1310_ sky130_fd_sc_hd__o211a_1
X_4393_ u_muldiv.o_div\[6\] net331 net377 net320 _2015_ VSS VSS VCC VCC _0257_
+ sky130_fd_sc_hd__a32o_1
X_3344_ net305 u_wr_mux.i_reg_data2\[20\] net563 VSS VSS VCC VCC net291 sky130_fd_sc_hd__mux2_1
X_3275_ _1210_ VSS VSS VCC VCC net196 sky130_fd_sc_hd__inv_4
X_5014_ clknet_leaf_35_i_clk _0047_ VSS VSS VCC VCC u_bits.i_op2\[3\] sky130_fd_sc_hd__dfxtp_1
X_4729_ net469 _2275_ _2278_ net488 VSS VSS VCC VCC _2279_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_143_i_clk clknet_4_8__leaf_i_clk VSS VSS VCC VCC clknet_leaf_143_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_158_i_clk clknet_4_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_158_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3060_ net574 _1023_ VSS VSS VCC VCC _1024_ sky130_fd_sc_hd__nor2_4
X_3962_ net307 net172 net388 VSS VSS VCC VCC _0124_ sky130_fd_sc_hd__mux2_1
X_2913_ _0468_ _0829_ _0471_ _0827_ VSS VSS VCC VCC _0884_ sky130_fd_sc_hd__a31o_1
X_3893_ net505 net96 net719 VSS VSS VCC VCC _1702_ sky130_fd_sc_hd__a21o_1
X_2844_ u_bits.i_op1\[22\] u_bits.i_op2\[22\] net411 _0786_ _0817_ vssd1 vssd1 vccd1
+ vccd1 _0818_ sky130_fd_sc_hd__a311o_1
X_2775_ _0749_ _0745_ _0489_ VSS VSS VCC VCC _0750_ sky130_fd_sc_hd__o21ai_2
X_4514_ u_muldiv.quotient_msk\[2\] net496 net342 u_muldiv.quotient_msk\[3\] vssd1
+ vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__a22o_1
X_4445_ net324 net375 _2051_ _2056_ VSS VSS VCC VCC _2057_ sky130_fd_sc_hd__o2bb2a_1
Xfanout604 net606 VSS VSS VCC VCC net604 sky130_fd_sc_hd__buf_4
X_4376_ u_muldiv.o_div\[3\] _1999_ net473 net496 VSS VSS VCC VCC _2002_ sky130_fd_sc_hd__o2bb2a_1
Xfanout615 net618 VSS VSS VCC VCC net615 sky130_fd_sc_hd__buf_2
Xfanout626 net633 VSS VSS VCC VCC net626 sky130_fd_sc_hd__buf_2
Xfanout637 net639 VSS VSS VCC VCC net637 sky130_fd_sc_hd__clkbuf_8
X_3327_ net39 _1254_ VSS VSS VCC VCC _0002_ sky130_fd_sc_hd__nor2_1
Xfanout648 net649 VSS VSS VCC VCC net648 sky130_fd_sc_hd__clkbuf_16
Xfanout659 u_bits.i_op1\[27\] VSS VSS VCC VCC net659 sky130_fd_sc_hd__clkbuf_8
X_3258_ _1198_ VSS VSS VCC VCC net186 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_60_i_clk clknet_4_7__leaf_i_clk VSS VSS VCC VCC clknet_leaf_60_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3189_ _1144_ _0907_ _0860_ net616 _1143_ VSS VSS VCC VCC _1145_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_75_i_clk clknet_4_13__leaf_i_clk VSS VSS VCC VCC clknet_leaf_75_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_13_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_13_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_28_i_clk clknet_4_4__leaf_i_clk VSS VSS VCC VCC clknet_leaf_28_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2560_ net448 net714 VSS VSS VCC VCC _0535_ sky130_fd_sc_hd__and2_1
Xoutput207 net207 VSS VSS VCC VCC o_add[31] sky130_fd_sc_hd__buf_2
Xoutput218 net218 VSS VSS VCC VCC o_instr_jal_jalr_branch sky130_fd_sc_hd__buf_2
Xoutput229 net229 VSS VSS VCC VCC o_pc_target[4] sky130_fd_sc_hd__buf_2
X_2491_ net446 u_bits.i_op2\[22\] VSS VSS VCC VCC _0466_ sky130_fd_sc_hd__and2_1
X_4230_ _0418_ net464 VSS VSS VCC VCC _1858_ sky130_fd_sc_hd__nand2_2
X_4161_ _0751_ _0752_ _1256_ VSS VSS VCC VCC _0205_ sky130_fd_sc_hd__and3_1
X_3112_ _1071_ _1072_ VSS VSS VCC VCC _1073_ sky130_fd_sc_hd__nand2_2
X_4092_ _1794_ u_bits.i_op2\[20\] _1787_ net380 VSS VSS VCC VCC _1800_ sky130_fd_sc_hd__o31a_1
X_3043_ u_bits.i_op2\[4\] _1006_ net328 VSS VSS VCC VCC _1007_ sky130_fd_sc_hd__o21a_1
X_4994_ clknet_leaf_48_i_clk _0027_ VSS VSS VCC VCC u_bits.i_op1\[24\] sky130_fd_sc_hd__dfxtp_1
X_3945_ net225 net129 net397 VSS VSS VCC VCC _0108_ sky130_fd_sc_hd__mux2_1
X_3876_ net507 _1688_ VSS VSS VCC VCC _1689_ sky130_fd_sc_hd__and2b_1
X_2827_ _0439_ _0438_ net645 VSS VSS VCC VCC _0801_ sky130_fd_sc_hd__mux2_1
X_2758_ _0724_ _0712_ _0725_ VSS VSS VCC VCC _0733_ sky130_fd_sc_hd__a21bo_1
X_2689_ net448 u_bits.i_op2\[15\] VSS VSS VCC VCC _0664_ sky130_fd_sc_hd__nand2_1
X_4428_ net436 _2042_ VSS VSS VCC VCC _2043_ sky130_fd_sc_hd__or2_1
Xfanout401 net402 VSS VSS VCC VCC net401 sky130_fd_sc_hd__buf_4
Xfanout412 _0782_ VSS VSS VCC VCC net412 sky130_fd_sc_hd__buf_6
Xfanout423 net426 VSS VSS VCC VCC net423 sky130_fd_sc_hd__buf_6
Xfanout434 net439 VSS VSS VCC VCC net434 sky130_fd_sc_hd__buf_6
Xfanout445 net446 VSS VSS VCC VCC net445 sky130_fd_sc_hd__buf_4
X_4359_ _1976_ _1977_ _1978_ _1986_ net329 VSS VSS VCC VCC _1987_ sky130_fd_sc_hd__o41ai_4
Xfanout456 net457 VSS VSS VCC VCC net456 sky130_fd_sc_hd__buf_4
Xfanout467 net468 VSS VSS VCC VCC net467 sky130_fd_sc_hd__buf_6
Xfanout478 net479 VSS VSS VCC VCC net478 sky130_fd_sc_hd__clkbuf_4
Xfanout489 net495 VSS VSS VCC VCC net489 sky130_fd_sc_hd__clkbuf_4
X_3730_ net578 _1606_ VSS VSS VCC VCC _1607_ sky130_fd_sc_hd__nor2_1
X_3661_ net530 _1533_ _1534_ _1542_ VSS VSS VCC VCC _1543_ sky130_fd_sc_hd__a31o_1
X_2612_ _0585_ _0586_ net429 VSS VSS VCC VCC _0587_ sky130_fd_sc_hd__a21oi_2
X_3592_ _1478_ u_pc_sel.i_pc_next\[11\] net575 VSS VSS VCC VCC net247 sky130_fd_sc_hd__mux2_8
X_5331_ clknet_leaf_143_i_clk _0359_ VSS VSS VCC VCC u_muldiv.divisor\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_2543_ _0517_ _0516_ _0515_ VSS VSS VCC VCC _0518_ sky130_fd_sc_hd__nand3b_1
X_5262_ clknet_leaf_119_i_clk _0290_ VSS VSS VCC VCC u_muldiv.quotient_msk\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2474_ u_muldiv.dividend\[25\] VSS VSS VCC VCC _0449_ sky130_fd_sc_hd__inv_2
X_4213_ op_cnt\[3\] op_cnt\[4\] op_cnt\[5\] _1838_ net510 VSS VSS VCC VCC
+ _1842_ sky130_fd_sc_hd__a41o_1
X_5193_ clknet_leaf_110_i_clk _0225_ VSS VSS VCC VCC u_muldiv.mul\[10\] sky130_fd_sc_hd__dfxtp_1
X_4144_ _1167_ _1168_ net406 VSS VSS VCC VCC _0188_ sky130_fd_sc_hd__a21oi_1
X_4075_ u_muldiv.divisor\[48\] net485 net336 u_muldiv.divisor\[49\] _1786_ vssd1 vssd1
+ vccd1 vccd1 _0168_ sky130_fd_sc_hd__a221o_1
X_3026_ net445 u_bits.i_op2\[27\] VSS VSS VCC VCC _0991_ sky130_fd_sc_hd__and2_1
X_4977_ clknet_leaf_47_i_clk _0010_ VSS VSS VCC VCC u_bits.i_op1\[7\] sky130_fd_sc_hd__dfxtp_4
X_3928_ net507 net574 net726 _1715_ VSS VSS VCC VCC _0092_ sky130_fd_sc_hd__o211a_4
X_3859_ u_bits.i_op2\[20\] net588 net548 VSS VSS VCC VCC _1676_ sky130_fd_sc_hd__mux2_1
X_4900_ u_muldiv.divisor\[7\] net492 net339 u_muldiv.divisor\[8\] vssd1 vssd1 vccd1
+ vccd1 _0352_ sky130_fd_sc_hd__a22o_1
X_4831_ u_muldiv.dividend\[26\] u_muldiv.dividend\[25\] u_muldiv.dividend\[24\] _2342_
+ VSS VSS VCC VCC _2372_ sky130_fd_sc_hd__or4_2
X_4762_ net679 net677 _2290_ net371 VSS VSS VCC VCC _2309_ sky130_fd_sc_hd__o31a_1
X_3713_ _1586_ _1590_ net520 VSS VSS VCC VCC _1591_ sky130_fd_sc_hd__a21oi_1
X_4693_ _1901_ _1902_ net459 VSS VSS VCC VCC _2246_ sky130_fd_sc_hd__a21o_1
X_3644_ _1526_ _1525_ net354 net189 VSS VSS VCC VCC _1527_ sky130_fd_sc_hd__a2bb2o_1
X_3575_ net443 _1459_ _1462_ net734 VSS VSS VCC VCC _1463_ sky130_fd_sc_hd__a211o_1
X_5314_ clknet_4_0__leaf_i_clk _0342_ VSS VSS VCC VCC u_muldiv.dividend\[29\]
+ sky130_fd_sc_hd__dfxtp_4
X_2526_ net641 net552 net681 net534 net424 VSS VSS VCC VCC _0501_ sky130_fd_sc_hd__o2111ai_1
X_5245_ clknet_4_8__leaf_i_clk _0273_ VSS VSS VCC VCC u_muldiv.o_div\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_2457_ net499 VSS VSS VCC VCC _0432_ sky130_fd_sc_hd__inv_6
X_5176_ clknet_leaf_59_i_clk _0208_ VSS VSS VCC VCC u_muldiv.add_prev\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_4127_ net583 net582 u_bits.i_op2\[28\] _1816_ VSS VSS VCC VCC _1827_ sky130_fd_sc_hd__or4_2
X_4058_ u_bits.i_op2\[14\] _1771_ _1772_ VSS VSS VCC VCC _1773_ sky130_fd_sc_hd__o21ba_1
X_3009_ net612 _0974_ _0890_ VSS VSS VCC VCC _0975_ sky130_fd_sc_hd__o21a_1
Xclkbuf_4_10__f_i_clk clknet_2_2_0_i_clk VSS VSS VCC VCC clknet_4_10__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3360_ net562 u_wr_mux.i_reg_data2\[30\] net418 net307 VSS VSS VCC VCC _1264_
+ sky130_fd_sc_hd__a22o_2
X_3291_ _1221_ VSS VSS VCC VCC net191 sky130_fd_sc_hd__inv_2
X_5030_ clknet_leaf_52_i_clk _0063_ VSS VSS VCC VCC u_bits.i_op2\[19\] sky130_fd_sc_hd__dfxtp_1
X_4814_ _1947_ _2355_ net465 VSS VSS VCC VCC _2356_ sky130_fd_sc_hd__o21ai_1
X_4745_ _2293_ net437 net326 net377 _2285_ VSS VSS VCC VCC _2294_ sky130_fd_sc_hd__a221oi_1
X_4676_ net489 _2230_ _2223_ net321 VSS VSS VCC VCC _2231_ sky130_fd_sc_hd__o211a_1
X_3627_ _0434_ _0781_ _0910_ _1113_ _1510_ VSS VSS VCC VCC _1511_ sky130_fd_sc_hd__o221a_1
X_3558_ net441 u_muldiv.mul\[41\] net413 _1446_ VSS VSS VCC VCC _1447_ sky130_fd_sc_hd__a31o_1
X_2509_ net531 _0430_ net517 net523 _0482_ VSS VSS VCC VCC _0484_ sky130_fd_sc_hd__o221ai_4
X_3489_ _0765_ _1381_ VSS VSS VCC VCC _1382_ sky130_fd_sc_hd__nand2_1
Xinput107 i_op2[8] VSS VSS VCC VCC net107 sky130_fd_sc_hd__buf_4
Xinput118 i_pc_next[4] VSS VSS VCC VCC net118 sky130_fd_sc_hd__clkbuf_1
X_5228_ clknet_leaf_115_i_clk _0256_ VSS VSS VCC VCC u_muldiv.o_div\[5\] sky130_fd_sc_hd__dfxtp_2
Xinput129 i_pc_target[15] VSS VSS VCC VCC net129 sky130_fd_sc_hd__clkbuf_1
X_5159_ clknet_4_14__leaf_i_clk _0191_ VSS VSS VCC VCC u_muldiv.add_prev\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2860_ _0832_ VSS VSS VCC VCC net198 sky130_fd_sc_hd__inv_6
X_2791_ net565 net558 net572 VSS VSS VCC VCC _0765_ sky130_fd_sc_hd__and3b_4
X_4530_ u_muldiv.quotient_msk\[18\] net490 net338 u_muldiv.quotient_msk\[19\] vssd1
+ vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__a22o_1
X_4461_ u_muldiv.o_div\[20\] _2069_ net319 VSS VSS VCC VCC _0271_ sky130_fd_sc_hd__mux2_1
X_3412_ net632 net717 net520 net352 VSS VSS VCC VCC _1309_ sky130_fd_sc_hd__a211o_1
X_4392_ net473 u_muldiv.quotient_msk\[6\] net438 _2013_ _2014_ VSS VSS VCC VCC
+ _2015_ sky130_fd_sc_hd__a32o_1
X_3343_ net304 u_wr_mux.i_reg_data2\[19\] net562 VSS VSS VCC VCC net289 sky130_fd_sc_hd__mux2_1
X_3274_ _0746_ _1209_ VSS VSS VCC VCC _1210_ sky130_fd_sc_hd__xor2_4
X_5013_ clknet_leaf_13_i_clk _0046_ VSS VSS VCC VCC u_bits.i_op2\[2\] sky130_fd_sc_hd__dfxtp_4
X_2989_ net23 net729 VSS VSS VCC VCC _0957_ sky130_fd_sc_hd__nor2_2
X_4728_ net682 _2276_ _2277_ VSS VSS VCC VCC _2278_ sky130_fd_sc_hd__o21a_1
X_4659_ _2206_ _0437_ _2114_ VSS VSS VCC VCC _2215_ sky130_fd_sc_hd__a21o_1
X_3961_ net306 net171 net399 VSS VSS VCC VCC _0123_ sky130_fd_sc_hd__mux2_1
X_2912_ _0878_ _0489_ VSS VSS VCC VCC _0883_ sky130_fd_sc_hd__nor2_1
X_3892_ net503 _1700_ VSS VSS VCC VCC _1701_ sky130_fd_sc_hd__and2b_1
X_2843_ _0796_ _0813_ _0816_ _0780_ VSS VSS VCC VCC _0817_ sky130_fd_sc_hd__a31o_1
X_2774_ _0480_ _0481_ _0488_ _0747_ VSS VSS VCC VCC _0749_ sky130_fd_sc_hd__nand4_4
X_4513_ u_muldiv.quotient_msk\[1\] net497 net342 u_muldiv.quotient_msk\[2\] vssd1
+ vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__a22o_1
X_4444_ net436 u_muldiv.quotient_msk\[17\] VSS VSS VCC VCC _2056_ sky130_fd_sc_hd__and2_1
X_4375_ _1998_ _2000_ _2001_ u_muldiv.o_div\[2\] VSS VSS VCC VCC _0253_ sky130_fd_sc_hd__o22a_1
Xfanout605 net606 VSS VSS VCC VCC net605 sky130_fd_sc_hd__clkbuf_2
Xfanout616 net618 VSS VSS VCC VCC net616 sky130_fd_sc_hd__buf_4
Xfanout627 net631 VSS VSS VCC VCC net627 sky130_fd_sc_hd__buf_4
X_3326_ net514 net2 _0432_ _1161_ VSS VSS VCC VCC _1254_ sky130_fd_sc_hd__o2bb2a_1
Xfanout638 net639 VSS VSS VCC VCC net638 sky130_fd_sc_hd__buf_2
Xfanout649 u_bits.i_op2\[0\] VSS VSS VCC VCC net649 sky130_fd_sc_hd__buf_6
X_3257_ _1193_ _1197_ VSS VSS VCC VCC _1198_ sky130_fd_sc_hd__nand2_8
Xclkbuf_leaf_9_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_9_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3188_ net651 net652 net654 net657 net639 net636 VSS VSS VCC VCC _1144_ sky130_fd_sc_hd__mux4_1
Xoutput208 net208 VSS VSS VCC VCC o_add[3] sky130_fd_sc_hd__buf_2
Xoutput219 net219 VSS VSS VCC VCC o_pc_select sky130_fd_sc_hd__buf_2
X_2490_ _0459_ net423 net671 net531 VSS VSS VCC VCC _0465_ sky130_fd_sc_hd__and4_1
X_4160_ net551 net500 net196 VSS VSS VCC VCC _0204_ sky130_fd_sc_hd__o21a_1
X_3111_ _1030_ _1035_ _1069_ _1029_ VSS VSS VCC VCC _1072_ sky130_fd_sc_hd__o211ai_2
X_4091_ _1794_ _0430_ _0429_ _0428_ VSS VSS VCC VCC _1799_ sky130_fd_sc_hd__and4b_2
X_3042_ net616 _1005_ net347 VSS VSS VCC VCC _1006_ sky130_fd_sc_hd__o21a_1
X_4993_ clknet_leaf_59_i_clk _0026_ VSS VSS VCC VCC u_bits.i_op1\[23\] sky130_fd_sc_hd__dfxtp_1
X_3944_ net224 net128 net396 VSS VSS VCC VCC _0107_ sky130_fd_sc_hd__mux2_1
X_3875_ u_bits.i_op2\[24\] u_bits.i_op2\[22\] net547 VSS VSS VCC VCC _1688_
+ sky130_fd_sc_hd__mux2_1
X_2826_ net645 _0437_ _0799_ VSS VSS VCC VCC _0800_ sky130_fd_sc_hd__o21a_1
X_2757_ _0630_ _0605_ _0729_ _0635_ VSS VSS VCC VCC _0732_ sky130_fd_sc_hd__o211ai_4
X_2688_ net647 net552 net687 net535 net423 VSS VSS VCC VCC _0663_ sky130_fd_sc_hd__o2111ai_2
Xclkbuf_leaf_142_i_clk clknet_4_8__leaf_i_clk VSS VSS VCC VCC clknet_leaf_142_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4427_ u_muldiv.o_div\[13\] u_muldiv.o_div\[14\] _2035_ VSS VSS VCC VCC _2042_
+ sky130_fd_sc_hd__nor3_2
Xfanout402 _1256_ VSS VSS VCC VCC net402 sky130_fd_sc_hd__buf_6
Xfanout413 net414 VSS VSS VCC VCC net413 sky130_fd_sc_hd__clkbuf_4
Xfanout424 net426 VSS VSS VCC VCC net424 sky130_fd_sc_hd__clkbuf_4
X_4358_ _1981_ _1983_ _1985_ _1984_ VSS VSS VCC VCC _1986_ sky130_fd_sc_hd__or4b_2
Xfanout435 net436 VSS VSS VCC VCC net435 sky130_fd_sc_hd__buf_4
Xfanout446 _0423_ VSS VSS VCC VCC net446 sky130_fd_sc_hd__buf_6
Xfanout457 _0420_ VSS VSS VCC VCC net457 sky130_fd_sc_hd__buf_6
X_3309_ _1128_ _1132_ VSS VSS VCC VCC _1239_ sky130_fd_sc_hd__nand2_1
Xfanout468 u_muldiv.on_wait VSS VSS VCC VCC net468 sky130_fd_sc_hd__buf_6
Xfanout479 net487 VSS VSS VCC VCC net479 sky130_fd_sc_hd__clkbuf_2
X_4289_ net462 u_muldiv.divisor\[17\] VSS VSS VCC VCC _1917_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_157_i_clk clknet_4_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_157_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3660_ _1219_ net356 net522 _1541_ net447 VSS VSS VCC VCC _1542_ sky130_fd_sc_hd__o221a_2
X_2611_ net449 net609 VSS VSS VCC VCC _0586_ sky130_fd_sc_hd__nand2_1
X_3591_ _1477_ net8 net733 VSS VSS VCC VCC _1478_ sky130_fd_sc_hd__mux2_1
X_5330_ clknet_leaf_137_i_clk _0358_ VSS VSS VCC VCC u_muldiv.divisor\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_2542_ net683 u_muldiv.add_prev\[17\] net535 VSS VSS VCC VCC _0517_ sky130_fd_sc_hd__mux2_1
X_5261_ clknet_leaf_117_i_clk _0289_ VSS VSS VCC VCC u_muldiv.quotient_msk\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2473_ u_muldiv.dividend\[27\] VSS VSS VCC VCC _0448_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_8__f_i_clk clknet_2_2_0_i_clk VSS VSS VCC VCC clknet_4_8__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4212_ op_cnt\[0\] op_cnt\[4\] _1159_ _1840_ net510 VSS VSS VCC VCC _0250_
+ sky130_fd_sc_hd__a311oi_1
Xclkbuf_leaf_74_i_clk clknet_4_13__leaf_i_clk VSS VSS VCC VCC clknet_leaf_74_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5192_ clknet_leaf_110_i_clk _0224_ VSS VSS VCC VCC u_muldiv.mul\[9\] sky130_fd_sc_hd__dfxtp_1
X_4143_ _1166_ _1169_ net401 VSS VSS VCC VCC _0187_ sky130_fd_sc_hd__and3_1
X_4074_ net589 _1784_ _1785_ VSS VSS VCC VCC _1786_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_89_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_89_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3025_ net732 net24 _0990_ VSS VSS VCC VCC net263 sky130_fd_sc_hd__o21a_4
Xclkbuf_leaf_12_i_clk clknet_4_4__leaf_i_clk VSS VSS VCC VCC clknet_leaf_12_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4976_ clknet_leaf_11_i_clk _0009_ VSS VSS VCC VCC u_bits.i_op1\[6\] sky130_fd_sc_hd__dfxtp_4
X_3927_ net178 net503 VSS VSS VCC VCC _1715_ sky130_fd_sc_hd__nand2b_2
X_3858_ net588 net728 _1675_ _1674_ VSS VSS VCC VCC _0062_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_27_i_clk clknet_4_4__leaf_i_clk VSS VSS VCC VCC clknet_leaf_27_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2809_ net572 net421 VSS VSS VCC VCC _0783_ sky130_fd_sc_hd__nand2_1
X_3789_ net509 net88 net722 VSS VSS VCC VCC _1624_ sky130_fd_sc_hd__a21o_1
X_4830_ u_muldiv.dividend\[25\] _2345_ u_muldiv.dividend\[26\] VSS VSS VCC VCC
+ _2371_ sky130_fd_sc_hd__o21ai_1
X_4761_ _1925_ _1936_ _2307_ VSS VSS VCC VCC _2308_ sky130_fd_sc_hd__o21ai_1
X_3712_ u_bits.i_op2\[20\] net675 net410 _1587_ _1589_ VSS VSS VCC VCC _1590_
+ sky130_fd_sc_hd__a311oi_4
X_4692_ _1902_ _1901_ VSS VSS VCC VCC _2245_ sky130_fd_sc_hd__nor2_1
X_3643_ _1524_ _1523_ _1520_ net521 VSS VSS VCC VCC _1526_ sky130_fd_sc_hd__a31o_1
X_3574_ net559 u_muldiv.mul\[10\] net413 net528 _1461_ VSS VSS VCC VCC _1462_
+ sky130_fd_sc_hd__o311a_1
X_5313_ clknet_leaf_170_i_clk _0341_ VSS VSS VCC VCC u_muldiv.dividend\[28\]
+ sky130_fd_sc_hd__dfxtp_2
X_2525_ net446 net588 VSS VSS VCC VCC _0500_ sky130_fd_sc_hd__nand2_1
X_5244_ clknet_leaf_152_i_clk _0272_ VSS VSS VCC VCC u_muldiv.o_div\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_2456_ u_bits.i_op2\[21\] VSS VSS VCC VCC _0431_ sky130_fd_sc_hd__inv_2
X_5175_ clknet_4_6__leaf_i_clk _0207_ VSS VSS VCC VCC u_muldiv.add_prev\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_4126_ u_muldiv.divisor\[59\] net482 net337 u_muldiv.divisor\[60\] _1826_ vssd1 vssd1
+ vccd1 vccd1 _0179_ sky130_fd_sc_hd__a221o_1
X_4057_ u_bits.i_op2\[14\] _1771_ net486 net468 VSS VSS VCC VCC _1772_ sky130_fd_sc_hd__a211o_1
X_3008_ _0771_ _0776_ net622 VSS VSS VCC VCC _0974_ sky130_fd_sc_hd__mux2_1
X_4959_ _0889_ net400 VSS VSS VCC VCC _0403_ sky130_fd_sc_hd__nor2_4
X_3290_ _0529_ _1220_ VSS VSS VCC VCC _1221_ sky130_fd_sc_hd__xnor2_4
X_4813_ _1944_ _1946_ _1945_ VSS VSS VCC VCC _2355_ sky130_fd_sc_hd__a21boi_1
X_4744_ net469 _2291_ _2292_ _2287_ _2288_ VSS VSS VCC VCC _2293_ sky130_fd_sc_hd__o32a_1
X_4675_ _2229_ _2228_ _2226_ _2224_ VSS VSS VCC VCC _2230_ sky130_fd_sc_hd__a2bb2o_1
X_3626_ u_bits.i_op2\[14\] net689 _1509_ VSS VSS VCC VCC _1510_ sky130_fd_sc_hd__o21ai_1
X_3557_ u_muldiv.dividend\[9\] net420 net368 u_muldiv.o_div\[9\] net360 vssd1 vssd1
+ vccd1 vccd1 _1446_ sky130_fd_sc_hd__a221o_1
X_2508_ net531 _0430_ _0482_ VSS VSS VCC VCC _0483_ sky130_fd_sc_hd__o21ai_1
X_3488_ _1379_ _1380_ net605 VSS VSS VCC VCC _1381_ sky130_fd_sc_hd__mux2_2
Xinput108 i_op2[9] VSS VSS VCC VCC net108 sky130_fd_sc_hd__buf_6
X_5227_ clknet_leaf_115_i_clk _0255_ VSS VSS VCC VCC u_muldiv.o_div\[4\] sky130_fd_sc_hd__dfxtp_2
Xinput119 i_pc_next[5] VSS VSS VCC VCC net119 sky130_fd_sc_hd__dlymetal6s2s_1
X_2439_ u_muldiv.divisor\[14\] VSS VSS VCC VCC _0414_ sky130_fd_sc_hd__inv_2
X_5158_ clknet_leaf_85_i_clk _0190_ VSS VSS VCC VCC u_muldiv.add_prev\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4109_ net586 net585 _1806_ net379 VSS VSS VCC VCC _1813_ sky130_fd_sc_hd__o31a_1
X_5089_ clknet_4_0__leaf_i_clk _0122_ VSS VSS VCC VCC net305 sky130_fd_sc_hd__dfxtp_4
X_2790_ net562 net570 VSS VSS VCC VCC _0764_ sky130_fd_sc_hd__and2b_4
X_4460_ _2066_ _2067_ net489 _2068_ VSS VSS VCC VCC _2069_ sky130_fd_sc_hd__a31o_1
X_3411_ net354 net194 _1306_ net412 _1307_ VSS VSS VCC VCC _1308_ sky130_fd_sc_hd__a2111o_1
X_4391_ u_muldiv.o_div\[5\] _2006_ u_muldiv.o_div\[6\] VSS VSS VCC VCC _2014_
+ sky130_fd_sc_hd__o21ai_1
X_3342_ net301 u_wr_mux.i_reg_data2\[18\] net562 VSS VSS VCC VCC net288 sky130_fd_sc_hd__mux2_8
X_3273_ _0748_ _0745_ _0488_ VSS VSS VCC VCC _1209_ sky130_fd_sc_hd__o21ai_2
X_5012_ clknet_leaf_40_i_clk _0045_ VSS VSS VCC VCC u_bits.i_op2\[1\] sky130_fd_sc_hd__dfxtp_2
X_2988_ net527 _0929_ _0930_ _0955_ VSS VSS VCC VCC _0956_ sky130_fd_sc_hd__a31o_1
X_4727_ _2276_ net682 net469 VSS VSS VCC VCC _2277_ sky130_fd_sc_hd__a21oi_1
X_4658_ _1888_ _2212_ _2213_ VSS VSS VCC VCC _2214_ sky130_fd_sc_hd__a21o_1
Xinput90 i_op2[21] VSS VSS VCC VCC net90 sky130_fd_sc_hd__buf_4
X_3609_ _1078_ net602 VSS VSS VCC VCC _1494_ sky130_fd_sc_hd__nand2b_1
X_4589_ u_muldiv.dividend\[4\] _2137_ u_muldiv.dividend\[5\] VSS VSS VCC VCC
+ _2151_ sky130_fd_sc_hd__o21ai_1
X_3960_ net305 net170 net386 VSS VSS VCC VCC _0122_ sky130_fd_sc_hd__mux2_1
X_2911_ _0742_ _0731_ _0880_ VSS VSS VCC VCC _0882_ sky130_fd_sc_hd__o21bai_4
X_3891_ u_bits.i_op2\[28\] net583 net545 VSS VSS VCC VCC _1700_ sky130_fd_sc_hd__mux2_1
X_2842_ net614 _0805_ net409 VSS VSS VCC VCC _0816_ sky130_fd_sc_hd__a21oi_1
X_2773_ _0488_ _0747_ VSS VSS VCC VCC _0748_ sky130_fd_sc_hd__nand2_2
X_4512_ net497 u_muldiv.quotient_msk\[0\] net342 u_muldiv.quotient_msk\[1\] vssd1
+ vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__a22o_1
X_4443_ u_muldiv.o_div\[17\] _2051_ net470 net491 VSS VSS VCC VCC _2055_ sky130_fd_sc_hd__o2bb2a_1
X_4374_ net325 net376 _1999_ u_muldiv.quotient_msk\[2\] VSS VSS VCC VCC _2001_
+ sky130_fd_sc_hd__o2bb2a_1
Xfanout606 net610 VSS VSS VCC VCC net606 sky130_fd_sc_hd__clkbuf_4
Xfanout617 net618 VSS VSS VCC VCC net617 sky130_fd_sc_hd__buf_4
X_3325_ _0433_ net512 net39 net486 VSS VSS VCC VCC _0001_ sky130_fd_sc_hd__a211o_1
Xfanout628 net630 VSS VSS VCC VCC net628 sky130_fd_sc_hd__clkbuf_4
Xfanout639 net640 VSS VSS VCC VCC net639 sky130_fd_sc_hd__buf_4
X_3256_ _1192_ _0649_ VSS VSS VCC VCC _1197_ sky130_fd_sc_hd__nand2_2
X_3187_ net623 _1014_ net452 VSS VSS VCC VCC _1143_ sky130_fd_sc_hd__and3_1
Xoutput209 net209 VSS VSS VCC VCC o_add[4] sky130_fd_sc_hd__buf_2
X_3110_ _1067_ _1068_ _1070_ VSS VSS VCC VCC _1071_ sky130_fd_sc_hd__nand3_1
X_4090_ u_muldiv.divisor\[51\] net484 net336 u_muldiv.divisor\[52\] _1798_ vssd1 vssd1
+ vccd1 vccd1 _0171_ sky130_fd_sc_hd__a221o_1
X_3041_ _0836_ _0841_ net623 VSS VSS VCC VCC _1005_ sky130_fd_sc_hd__mux2_1
X_4992_ clknet_leaf_46_i_clk _0025_ VSS VSS VCC VCC u_bits.i_op1\[22\] sky130_fd_sc_hd__dfxtp_4
X_3943_ net223 net127 net397 VSS VSS VCC VCC _0106_ sky130_fd_sc_hd__mux2_1
X_3874_ u_bits.i_op2\[22\] net724 _1687_ _1686_ VSS VSS VCC VCC _0066_ sky130_fd_sc_hd__o22a_1
X_2825_ net645 net699 VSS VSS VCC VCC _0799_ sky130_fd_sc_hd__nand2_1
X_2756_ _0636_ _0637_ _0730_ VSS VSS VCC VCC _0731_ sky130_fd_sc_hd__a21oi_2
X_2687_ _0656_ _0659_ _0658_ _0646_ _0648_ VSS VSS VCC VCC _0662_ sky130_fd_sc_hd__o2111ai_4
X_4426_ net318 _2039_ _2041_ VSS VSS VCC VCC _0264_ sky130_fd_sc_hd__a21oi_1
Xfanout403 net408 VSS VSS VCC VCC net403 sky130_fd_sc_hd__buf_4
Xfanout414 net415 VSS VSS VCC VCC net414 sky130_fd_sc_hd__buf_4
Xfanout425 net426 VSS VSS VCC VCC net425 sky130_fd_sc_hd__buf_12
X_4357_ u_muldiv.divisor\[47\] u_muldiv.divisor\[46\] u_muldiv.divisor\[45\] u_muldiv.divisor\[44\]
+ VSS VSS VCC VCC _1985_ sky130_fd_sc_hd__or4_2
Xfanout436 net439 VSS VSS VCC VCC net436 sky130_fd_sc_hd__buf_4
Xfanout447 net449 VSS VSS VCC VCC net447 sky130_fd_sc_hd__buf_4
X_3308_ _1138_ _1139_ _1237_ VSS VSS VCC VCC _1238_ sky130_fd_sc_hd__nand3_1
Xfanout458 _0419_ VSS VSS VCC VCC net458 sky130_fd_sc_hd__buf_6
X_4288_ u_muldiv.divisor\[17\] net462 VSS VSS VCC VCC _1916_ sky130_fd_sc_hd__nand2b_1
Xfanout469 net472 VSS VSS VCC VCC net469 sky130_fd_sc_hd__buf_4
X_3239_ _1183_ VSS VSS VCC VCC net213 sky130_fd_sc_hd__clkinv_8
X_2610_ net648 net554 net710 net539 net425 VSS VSS VCC VCC _0585_ sky130_fd_sc_hd__o2111ai_2
Xclkbuf_leaf_8_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_8_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3590_ net530 _1473_ _1475_ _1476_ VSS VSS VCC VCC _1477_ sky130_fd_sc_hd__a2bb2o_1
X_2541_ _0511_ _0512_ net432 VSS VSS VCC VCC _0516_ sky130_fd_sc_hd__o21ai_1
X_5260_ clknet_leaf_116_i_clk _0288_ VSS VSS VCC VCC u_muldiv.quotient_msk\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2472_ u_muldiv.dividend\[30\] VSS VSS VCC VCC _0447_ sky130_fd_sc_hd__inv_2
X_4211_ op_cnt\[3\] op_cnt\[4\] _1838_ VSS VSS VCC VCC _1841_ sky130_fd_sc_hd__and3_1
X_5191_ clknet_4_11__leaf_i_clk _0223_ VSS VSS VCC VCC u_muldiv.mul\[8\] sky130_fd_sc_hd__dfxtp_1
X_4142_ _1162_ _1163_ net406 VSS VSS VCC VCC _0186_ sky130_fd_sc_hd__a21oi_1
X_4073_ net589 _1784_ net384 VSS VSS VCC VCC _1785_ sky130_fd_sc_hd__o21ai_1
X_3024_ net735 _0989_ net574 VSS VSS VCC VCC _0990_ sky130_fd_sc_hd__o21ba_4
X_4975_ clknet_leaf_43_i_clk _0008_ VSS VSS VCC VCC u_bits.i_op1\[5\] sky130_fd_sc_hd__dfxtp_4
X_3926_ net502 net242 net723 _1714_ VSS VSS VCC VCC _0091_ sky130_fd_sc_hd__o211a_1
X_3857_ net513 net86 net721 VSS VSS VCC VCC _1675_ sky130_fd_sc_hd__a21o_1
X_2808_ net566 net558 net572 VSS VSS VCC VCC _0782_ sky130_fd_sc_hd__and3_4
X_3788_ net509 _1622_ VSS VSS VCC VCC _1623_ sky130_fd_sc_hd__and2b_1
X_2739_ _0711_ _0710_ _0709_ VSS VSS VCC VCC _0714_ sky130_fd_sc_hd__nand3b_2
X_4409_ u_muldiv.o_div\[9\] u_muldiv.o_div\[10\] _2020_ net492 VSS VSS VCC VCC
+ _2028_ sky130_fd_sc_hd__o31a_1
X_4760_ _1925_ _1936_ net459 VSS VSS VCC VCC _2307_ sky130_fd_sc_hd__a21oi_1
X_3711_ u_bits.i_op2\[20\] net676 net349 _1588_ VSS VSS VCC VCC _1589_ sky130_fd_sc_hd__o211a_2
X_4691_ _2242_ _2243_ net489 VSS VSS VCC VCC _2244_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_156_i_clk clknet_4_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_156_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3642_ u_bits.i_op2\[15\] net687 net352 VSS VSS VCC VCC _1525_ sky130_fd_sc_hd__a21oi_1
X_3573_ u_muldiv.o_div\[10\] net366 net358 _1460_ VSS VSS VCC VCC _1461_ sky130_fd_sc_hd__a211o_1
X_5312_ clknet_leaf_170_i_clk _0340_ VSS VSS VCC VCC u_muldiv.dividend\[27\]
+ sky130_fd_sc_hd__dfxtp_2
X_2524_ _0497_ _0498_ VSS VSS VCC VCC _0499_ sky130_fd_sc_hd__nand2_2
X_2455_ u_bits.i_op2\[20\] VSS VSS VCC VCC _0430_ sky130_fd_sc_hd__inv_2
X_5243_ clknet_leaf_153_i_clk _0271_ VSS VSS VCC VCC u_muldiv.o_div\[20\]
+ sky130_fd_sc_hd__dfxtp_2
X_5174_ clknet_4_6__leaf_i_clk _0206_ VSS VSS VCC VCC u_muldiv.add_prev\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_4125_ u_bits.i_op2\[28\] _1824_ _1825_ VSS VSS VCC VCC _1826_ sky130_fd_sc_hd__a21oi_1
X_4056_ net593 net592 _1764_ net381 VSS VSS VCC VCC _1771_ sky130_fd_sc_hd__o31a_1
X_3007_ net522 _0760_ net201 VSS VSS VCC VCC _0973_ sky130_fd_sc_hd__o21a_1
X_4958_ _1256_ _0832_ VSS VSS VCC VCC _0402_ sky130_fd_sc_hd__nor2_4
X_3909_ net579 net720 _1712_ _1713_ VSS VSS VCC VCC _0075_ sky130_fd_sc_hd__a211o_1
X_4889_ u_muldiv.dividend\[30\] _2402_ u_muldiv.dividend\[31\] VSS VSS VCC VCC
+ _2425_ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_73_i_clk clknet_4_13__leaf_i_clk VSS VSS VCC VCC clknet_leaf_73_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_11_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_11_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_26_i_clk clknet_4_6__leaf_i_clk VSS VSS VCC VCC clknet_leaf_26_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4812_ u_muldiv.dividend\[24\] _2354_ _1993_ VSS VSS VCC VCC _0337_ sky130_fd_sc_hd__mux2_1
X_4743_ _2290_ net371 net679 VSS VSS VCC VCC _2292_ sky130_fd_sc_hd__a21oi_1
X_4674_ _2227_ net372 net693 net469 VSS VSS VCC VCC _2229_ sky130_fd_sc_hd__a31o_1
X_3625_ net564 _1508_ net350 VSS VSS VCC VCC _1509_ sky130_fd_sc_hd__o21a_1
X_3556_ _1181_ net356 net521 _1444_ VSS VSS VCC VCC _1445_ sky130_fd_sc_hd__o22a_2
X_2507_ net646 net553 net676 net531 net423 VSS VSS VCC VCC _0482_ sky130_fd_sc_hd__o2111ai_4
X_3487_ _0767_ _0931_ _0932_ _1294_ net453 net450 VSS VSS VCC VCC _1380_ sky130_fd_sc_hd__mux4_2
X_5226_ clknet_leaf_96_i_clk _0254_ VSS VSS VCC VCC u_muldiv.o_div\[3\] sky130_fd_sc_hd__dfxtp_1
Xinput109 i_pc_next[10] VSS VSS VCC VCC net109 sky130_fd_sc_hd__clkbuf_1
X_2438_ net470 VSS VSS VCC VCC _0413_ sky130_fd_sc_hd__clkinv_4
X_5157_ clknet_leaf_86_i_clk _0189_ VSS VSS VCC VCC u_muldiv.add_prev\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4108_ u_muldiv.divisor\[55\] net439 _1720_ u_muldiv.divisor\[56\] _1812_ vssd1 vssd1
+ vccd1 vccd1 _0175_ sky130_fd_sc_hd__o221a_1
X_5088_ clknet_leaf_11_i_clk _0121_ VSS VSS VCC VCC net304 sky130_fd_sc_hd__dfxtp_4
X_4039_ net595 _1757_ net484 net468 VSS VSS VCC VCC _1758_ sky130_fd_sc_hd__a211o_1
X_3410_ net572 net368 _1303_ _1304_ VSS VSS VCC VCC _1307_ sky130_fd_sc_hd__a31o_1
X_4390_ u_muldiv.o_div\[5\] u_muldiv.o_div\[6\] _2006_ net493 VSS VSS VCC VCC
+ _2013_ sky130_fd_sc_hd__o31a_1
X_3341_ net290 u_wr_mux.i_reg_data2\[17\] net562 VSS VSS VCC VCC net287 sky130_fd_sc_hd__mux2_4
X_3272_ _0509_ _1206_ VSS VSS VCC VCC net192 sky130_fd_sc_hd__xor2_4
X_5011_ clknet_leaf_15_i_clk _0044_ VSS VSS VCC VCC u_bits.i_op2\[0\] sky130_fd_sc_hd__dfxtp_4
X_2987_ net522 _0954_ net356 _0928_ net442 VSS VSS VCC VCC _0955_ sky130_fd_sc_hd__o221a_1
X_4726_ net684 _2267_ net373 VSS VSS VCC VCC _2276_ sky130_fd_sc_hd__o21ai_1
X_4657_ _1888_ _2212_ net470 VSS VSS VCC VCC _2213_ sky130_fd_sc_hd__o21ai_1
Xinput80 i_op2[12] VSS VSS VCC VCC net80 sky130_fd_sc_hd__dlymetal6s2s_1
X_3608_ net592 net691 _1492_ net348 VSS VSS VCC VCC _1493_ sky130_fd_sc_hd__o211a_1
Xinput91 i_op2[22] VSS VSS VCC VCC net91 sky130_fd_sc_hd__buf_2
X_4588_ u_muldiv.dividend\[3\] u_muldiv.dividend\[5\] u_muldiv.dividend\[4\] _2126_
+ VSS VSS VCC VCC _2150_ sky130_fd_sc_hd__or4_1
X_3539_ _1428_ _1426_ _0910_ _0900_ VSS VSS VCC VCC _1429_ sky130_fd_sc_hd__o2bb2a_2
X_5209_ clknet_leaf_156_i_clk _0241_ VSS VSS VCC VCC u_muldiv.mul\[26\] sky130_fd_sc_hd__dfxtp_1
X_2910_ _0880_ VSS VSS VCC VCC _0881_ sky130_fd_sc_hd__inv_2
X_3890_ net583 net723 _1699_ _1698_ VSS VSS VCC VCC _0070_ sky130_fd_sc_hd__o22a_1
X_2841_ net564 net558 net573 VSS VSS VCC VCC _0815_ sky130_fd_sc_hd__or3b_2
X_2772_ _0484_ _0485_ _0487_ VSS VSS VCC VCC _0747_ sky130_fd_sc_hd__nand3_2
X_4511_ net323 _2106_ _2108_ VSS VSS VCC VCC _0282_ sky130_fd_sc_hd__o21a_1
X_4442_ u_muldiv.o_div\[16\] net324 net375 _2054_ VSS VSS VCC VCC _0267_ sky130_fd_sc_hd__a31o_1
X_4373_ u_muldiv.o_div\[2\] _1994_ _1999_ VSS VSS VCC VCC _2000_ sky130_fd_sc_hd__a21boi_1
Xfanout607 net610 VSS VSS VCC VCC net607 sky130_fd_sc_hd__clkbuf_4
Xfanout618 u_bits.i_op2\[3\] VSS VSS VCC VCC net618 sky130_fd_sc_hd__buf_8
X_3324_ net39 _1253_ VSS VSS VCC VCC net219 sky130_fd_sc_hd__nor2_4
Xfanout629 net630 VSS VSS VCC VCC net629 sky130_fd_sc_hd__buf_2
X_3255_ _1196_ VSS VSS VCC VCC net187 sky130_fd_sc_hd__inv_2
X_3186_ u_muldiv.mul\[63\] net363 net357 u_muldiv.mul\[31\] _1141_ vssd1 vssd1 vccd1
+ vccd1 _1142_ sky130_fd_sc_hd__a221o_1
X_4709_ u_muldiv.dividend\[15\] _2260_ net319 VSS VSS VCC VCC _0328_ sky130_fd_sc_hd__mux2_1
X_3040_ u_muldiv.mul\[59\] net363 net357 u_muldiv.mul\[27\] _1003_ vssd1 vssd1 vccd1
+ vccd1 _1004_ sky130_fd_sc_hd__a221o_1
X_4991_ clknet_leaf_137_i_clk _0024_ VSS VSS VCC VCC u_bits.i_op1\[21\] sky130_fd_sc_hd__dfxtp_1
X_3942_ net222 net126 net393 VSS VSS VCC VCC _0105_ sky130_fd_sc_hd__mux2_1
X_3873_ net502 net91 net720 VSS VSS VCC VCC _1687_ sky130_fd_sc_hd__a21o_1
X_2824_ net458 net701 _0797_ VSS VSS VCC VCC _0798_ sky130_fd_sc_hd__a21oi_1
X_2755_ _0685_ _0728_ VSS VSS VCC VCC _0730_ sky130_fd_sc_hd__nand2_1
X_2686_ _0660_ VSS VSS VCC VCC _0661_ sky130_fd_sc_hd__inv_2
X_4425_ net318 _2040_ u_muldiv.o_div\[13\] VSS VSS VCC VCC _2041_ sky130_fd_sc_hd__a21oi_1
Xfanout404 net408 VSS VSS VCC VCC net404 sky130_fd_sc_hd__buf_6
X_4356_ u_muldiv.dividend\[31\] u_muldiv.divisor\[31\] VSS VSS VCC VCC _1984_
+ sky130_fd_sc_hd__nand2b_2
Xfanout415 _0758_ VSS VSS VCC VCC net415 sky130_fd_sc_hd__buf_2
Xfanout426 _0461_ VSS VSS VCC VCC net426 sky130_fd_sc_hd__clkbuf_8
Xfanout437 net439 VSS VSS VCC VCC net437 sky130_fd_sc_hd__buf_4
Xfanout448 net449 VSS VSS VCC VCC net448 sky130_fd_sc_hd__buf_4
X_3307_ _1128_ _1132_ VSS VSS VCC VCC _1237_ sky130_fd_sc_hd__or2_1
Xfanout459 _0413_ VSS VSS VCC VCC net459 sky130_fd_sc_hd__buf_12
X_4287_ _1913_ _1914_ VSS VSS VCC VCC _1915_ sky130_fd_sc_hd__nor2_1
X_3238_ _1178_ _1182_ VSS VSS VCC VCC _1183_ sky130_fd_sc_hd__nand2b_4
X_3169_ _1126_ net29 net733 VSS VSS VCC VCC _1127_ sky130_fd_sc_hd__mux2_1
X_2540_ net535 net683 _0463_ _0511_ net432 VSS VSS VCC VCC _0515_ sky130_fd_sc_hd__a311o_1
X_2471_ u_muldiv.dividend\[10\] VSS VSS VCC VCC _0446_ sky130_fd_sc_hd__inv_2
X_4210_ op_cnt\[3\] _1838_ op_cnt\[4\] VSS VSS VCC VCC _1840_ sky130_fd_sc_hd__a21oi_1
X_5190_ clknet_leaf_112_i_clk _0222_ VSS VSS VCC VCC u_muldiv.mul\[7\] sky130_fd_sc_hd__dfxtp_1
X_4141_ net555 net500 net205 VSS VSS VCC VCC _0185_ sky130_fd_sc_hd__o21a_1
X_4072_ net591 net590 _1775_ net380 VSS VSS VCC VCC _1784_ sky130_fd_sc_hd__o31a_1
X_3023_ net544 _0973_ _0988_ _0972_ VSS VSS VCC VCC _0989_ sky130_fd_sc_hd__o31a_1
X_4974_ clknet_leaf_90_i_clk _0007_ VSS VSS VCC VCC u_bits.i_op1\[4\] sky130_fd_sc_hd__dfxtp_2
X_3925_ net177 net504 VSS VSS VCC VCC _1714_ sky130_fd_sc_hd__nand2b_1
X_3856_ net512 _1673_ VSS VSS VCC VCC _1674_ sky130_fd_sc_hd__and2b_1
X_2807_ net560 net570 VSS VSS VCC VCC _0781_ sky130_fd_sc_hd__nand2_8
X_3787_ net624 net641 net548 VSS VSS VCC VCC _1622_ sky130_fd_sc_hd__mux2_1
X_2738_ _0709_ _0710_ _0711_ VSS VSS VCC VCC _0713_ sky130_fd_sc_hd__a21bo_1
X_2669_ _0640_ _0641_ net519 net526 VSS VSS VCC VCC _0644_ sky130_fd_sc_hd__a211o_1
X_4408_ u_muldiv.o_div\[7\] _0452_ _2012_ _0453_ VSS VSS VCC VCC _2027_ sky130_fd_sc_hd__and4b_1
X_4339_ _1961_ _1966_ _1963_ VSS VSS VCC VCC _1967_ sky130_fd_sc_hd__or3b_1
X_3710_ _0430_ net569 net676 VSS VSS VCC VCC _1588_ sky130_fd_sc_hd__or3b_1
X_4690_ u_muldiv.dividend\[13\] u_muldiv.dividend\[12\] _2218_ u_muldiv.dividend\[14\]
+ VSS VSS VCC VCC _2243_ sky130_fd_sc_hd__o31a_1
X_3641_ net608 net409 _1150_ net440 _0781_ VSS VSS VCC VCC _1524_ sky130_fd_sc_hd__o32a_1
X_3572_ net567 net556 u_muldiv.dividend\[10\] u_muldiv.mul\[42\] net362 vssd1 vssd1
+ vccd1 vccd1 _1460_ sky130_fd_sc_hd__a32o_1
X_5311_ clknet_leaf_170_i_clk _0339_ VSS VSS VCC VCC u_muldiv.dividend\[26\]
+ sky130_fd_sc_hd__dfxtp_2
X_2523_ _0492_ _0493_ _0495_ VSS VSS VCC VCC _0498_ sky130_fd_sc_hd__nand3_2
X_5242_ clknet_leaf_139_i_clk _0270_ VSS VSS VCC VCC u_muldiv.o_div\[19\]
+ sky130_fd_sc_hd__dfxtp_2
X_2454_ net589 VSS VSS VCC VCC _0429_ sky130_fd_sc_hd__inv_2
X_5173_ clknet_leaf_70_i_clk _0205_ VSS VSS VCC VCC u_muldiv.add_prev\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_4124_ u_bits.i_op2\[28\] _1824_ net384 VSS VSS VCC VCC _1825_ sky130_fd_sc_hd__o21ai_1
Xinput1 i_alu_ctrl[0] VSS VSS VCC VCC net1 sky130_fd_sc_hd__clkbuf_1
X_4055_ u_muldiv.divisor\[44\] net485 net335 u_muldiv.divisor\[45\] _1770_ vssd1 vssd1
+ vccd1 vccd1 _0164_ sky130_fd_sc_hd__a221o_1
X_3006_ u_muldiv.mul\[58\] net363 net357 u_muldiv.mul\[26\] _0971_ vssd1 vssd1 vccd1
+ vccd1 _0972_ sky130_fd_sc_hd__a221o_1
X_4957_ _0751_ _0752_ net407 VSS VSS VCC VCC _0401_ sky130_fd_sc_hd__and3_1
X_3908_ net501 net580 net545 net723 VSS VSS VCC VCC _1713_ sky130_fd_sc_hd__and4b_1
X_4888_ _2419_ _2421_ net466 _2423_ net479 VSS VSS VCC VCC _2424_ sky130_fd_sc_hd__a311oi_1
X_3839_ net591 net592 net547 VSS VSS VCC VCC _1661_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_7_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_7_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4811_ net480 _2345_ _2346_ _2353_ VSS VSS VCC VCC _2354_ sky130_fd_sc_hd__a31o_1
X_4742_ net684 net682 _2267_ net373 net679 VSS VSS VCC VCC _2291_ sky130_fd_sc_hd__o311a_1
X_4673_ _2227_ net372 net693 VSS VSS VCC VCC _2228_ sky130_fd_sc_hd__a21oi_1
X_3624_ u_bits.i_op2\[14\] net689 VSS VSS VCC VCC _1508_ sky130_fd_sc_hd__nand2_1
X_3555_ net353 _1440_ _1442_ _1443_ VSS VSS VCC VCC _1444_ sky130_fd_sc_hd__a31o_1
X_2506_ _0477_ _0478_ _0479_ VSS VSS VCC VCC _0481_ sky130_fd_sc_hd__a21o_1
X_3486_ _1293_ _1297_ _1298_ _1301_ net453 net450 VSS VSS VCC VCC _1379_ sky130_fd_sc_hd__mux4_1
X_5225_ clknet_leaf_95_i_clk _0253_ VSS VSS VCC VCC u_muldiv.o_div\[2\] sky130_fd_sc_hd__dfxtp_2
X_5156_ clknet_leaf_102_i_clk _0188_ VSS VSS VCC VCC u_muldiv.add_prev\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4107_ net585 _1810_ _1811_ VSS VSS VCC VCC _1812_ sky130_fd_sc_hd__a21o_1
X_5087_ clknet_leaf_34_i_clk _0120_ VSS VSS VCC VCC net301 sky130_fd_sc_hd__dfxtp_4
X_4038_ net597 net596 _1749_ net379 VSS VSS VCC VCC _1757_ sky130_fd_sc_hd__o31a_1
Xoutput190 net190 VSS VSS VCC VCC o_add[16] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_155_i_clk clknet_4_9__leaf_i_clk VSS VSS VCC VCC clknet_leaf_155_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3340_ net279 u_wr_mux.i_reg_data2\[16\] net565 VSS VSS VCC VCC net286 sky130_fd_sc_hd__mux2_4
X_3271_ _1208_ VSS VSS VCC VCC net193 sky130_fd_sc_hd__inv_2
X_5010_ clknet_leaf_24_i_clk _0043_ VSS VSS VCC VCC u_pc_sel.i_inst_branch
+ sky130_fd_sc_hd__dfxtp_1
X_2986_ _0901_ _0941_ _0949_ _0953_ VSS VSS VCC VCC _0954_ sky130_fd_sc_hd__o211a_1
X_4725_ _1917_ _2273_ _2274_ VSS VSS VCC VCC _2275_ sky130_fd_sc_hd__o21a_1
X_4656_ _1885_ _2203_ VSS VSS VCC VCC _2212_ sky130_fd_sc_hd__or2_1
Xinput70 i_op1[3] VSS VSS VCC VCC net70 sky130_fd_sc_hd__clkbuf_1
X_3607_ net564 net691 u_bits.i_op2\[13\] VSS VSS VCC VCC _1492_ sky130_fd_sc_hd__nand3b_1
Xinput81 i_op2[13] VSS VSS VCC VCC net81 sky130_fd_sc_hd__clkbuf_2
X_4587_ u_muldiv.dividend\[4\] _2149_ net320 VSS VSS VCC VCC _0317_ sky130_fd_sc_hd__mux2_1
Xinput92 i_op2[23] VSS VSS VCC VCC net92 sky130_fd_sc_hd__buf_6
X_3538_ net604 _1427_ net365 net573 VSS VSS VCC VCC _1428_ sky130_fd_sc_hd__o211a_1
X_3469_ net453 _0891_ _1362_ VSS VSS VCC VCC _1363_ sky130_fd_sc_hd__o21ai_2
X_5208_ clknet_leaf_156_i_clk _0240_ VSS VSS VCC VCC u_muldiv.mul\[25\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_72_i_clk clknet_4_13__leaf_i_clk VSS VSS VCC VCC clknet_leaf_72_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5139_ clknet_leaf_42_i_clk _0171_ VSS VSS VCC VCC u_muldiv.divisor\[51\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_87_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_87_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_10_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_10_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2840_ net560 net440 net571 VSS VSS VCC VCC _0814_ sky130_fd_sc_hd__and3b_4
X_2771_ _0480_ _0481_ VSS VSS VCC VCC _0746_ sky130_fd_sc_hd__nand2_2
X_4510_ net315 _2107_ u_muldiv.o_div\[31\] VSS VSS VCC VCC _2108_ sky130_fd_sc_hd__a21o_1
X_4441_ net324 net375 _2052_ _2053_ VSS VSS VCC VCC _2054_ sky130_fd_sc_hd__o2bb2a_1
X_4372_ u_muldiv.o_div\[0\] u_muldiv.o_div\[1\] u_muldiv.o_div\[2\] net496 vssd1 vssd1
+ vccd1 vccd1 _1999_ sky130_fd_sc_hd__o31a_1
X_3323_ _1245_ _1252_ u_pc_sel.i_inst_branch u_pc_sel.i_inst_jal_jalr vssd1 vssd1
+ vccd1 vccd1 _1253_ sky130_fd_sc_hd__a31oi_4
Xfanout608 net609 VSS VSS VCC VCC net608 sky130_fd_sc_hd__clkbuf_4
Xfanout619 net622 VSS VSS VCC VCC net619 sky130_fd_sc_hd__clkbuf_4
X_3254_ _1194_ _1195_ VSS VSS VCC VCC _1196_ sky130_fd_sc_hd__nand2_4
X_3185_ u_muldiv.dividend\[31\] net419 net364 u_muldiv.o_div\[31\] net442 vssd1 vssd1
+ vccd1 vccd1 _1141_ sky130_fd_sc_hd__a221o_2
X_2969_ net708 net710 net713 net715 net643 net628 VSS VSS VCC VCC _0937_ sky130_fd_sc_hd__mux4_1
X_4708_ net488 _2258_ _2259_ _2257_ VSS VSS VCC VCC _2260_ sky130_fd_sc_hd__a31o_1
X_4639_ net699 _2195_ net385 VSS VSS VCC VCC _2197_ sky130_fd_sc_hd__o21ai_1
X_4990_ clknet_leaf_132_i_clk _0023_ VSS VSS VCC VCC u_bits.i_op1\[20\] sky130_fd_sc_hd__dfxtp_4
X_3941_ net221 net125 net397 VSS VSS VCC VCC _0104_ sky130_fd_sc_hd__mux2_1
X_3872_ net503 _1685_ VSS VSS VCC VCC _1686_ sky130_fd_sc_hd__and2b_1
X_2823_ net458 _0436_ VSS VSS VCC VCC _0797_ sky130_fd_sc_hd__nor2_1
X_2754_ _0662_ _0684_ _0706_ _0726_ VSS VSS VCC VCC _0729_ sky130_fd_sc_hd__nor4_4
X_2685_ _0656_ _0659_ _0658_ VSS VSS VCC VCC _0660_ sky130_fd_sc_hd__o21ai_4
X_4424_ _2035_ u_muldiv.quotient_msk\[13\] net436 VSS VSS VCC VCC _2040_ sky130_fd_sc_hd__mux2_1
X_4355_ _1979_ _1980_ _1982_ VSS VSS VCC VCC _1983_ sky130_fd_sc_hd__or3_1
Xfanout405 net408 VSS VSS VCC VCC net405 sky130_fd_sc_hd__buf_4
Xfanout416 net418 VSS VSS VCC VCC net416 sky130_fd_sc_hd__buf_12
Xfanout427 net430 VSS VSS VCC VCC net427 sky130_fd_sc_hd__buf_6
X_3306_ _1224_ _1235_ net440 VSS VSS VCC VCC _1236_ sky130_fd_sc_hd__o21a_1
Xfanout438 net439 VSS VSS VCC VCC net438 sky130_fd_sc_hd__buf_4
Xfanout449 _0423_ VSS VSS VCC VCC net449 sky130_fd_sc_hd__buf_4
X_4286_ u_muldiv.dividend\[16\] u_muldiv.divisor\[16\] VSS VSS VCC VCC _1914_
+ sky130_fd_sc_hd__and2b_1
X_3237_ _0636_ _0637_ _0715_ VSS VSS VCC VCC _1182_ sky130_fd_sc_hd__nand3_1
X_3168_ _1111_ _1112_ net527 _1125_ VSS VSS VCC VCC _1126_ sky130_fd_sc_hd__o22a_4
X_3099_ net735 _1060_ net575 VSS VSS VCC VCC _1061_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_4_13__f_i_clk clknet_2_3_0_i_clk VSS VSS VCC VCC clknet_4_13__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2470_ u_muldiv.dividend\[12\] VSS VSS VCC VCC _0445_ sky130_fd_sc_hd__clkinv_2
X_4140_ net555 net500 net194 VSS VSS VCC VCC _0184_ sky130_fd_sc_hd__o21a_1
X_4071_ u_muldiv.divisor\[47\] net485 net336 u_muldiv.divisor\[48\] _1783_ vssd1 vssd1
+ vccd1 vccd1 _0167_ sky130_fd_sc_hd__a221o_1
X_3022_ _0977_ _0985_ _0987_ _0422_ VSS VSS VCC VCC _0988_ sky130_fd_sc_hd__o31a_1
X_4973_ clknet_leaf_78_i_clk _0006_ VSS VSS VCC VCC u_bits.i_op1\[3\] sky130_fd_sc_hd__dfxtp_1
X_3924_ u_pc_sel.i_pc_next\[15\] net114 net389 VSS VSS VCC VCC _0090_ sky130_fd_sc_hd__mux2_1
X_3855_ u_bits.i_op2\[19\] net589 net548 VSS VSS VCC VCC _1673_ sky130_fd_sc_hd__mux2_1
X_2806_ net606 _0778_ net327 VSS VSS VCC VCC _0780_ sky130_fd_sc_hd__o21a_1
X_3786_ net640 net719 _1620_ _1621_ VSS VSS VCC VCC _0044_ sky130_fd_sc_hd__a211o_1
X_2737_ _0709_ _0710_ _0711_ VSS VSS VCC VCC _0712_ sky130_fd_sc_hd__a21boi_2
X_2668_ _0640_ _0641_ net432 VSS VSS VCC VCC _0643_ sky130_fd_sc_hd__a21o_1
X_4407_ net318 _2024_ _2026_ VSS VSS VCC VCC _0260_ sky130_fd_sc_hd__a21oi_1
X_2599_ net537 u_muldiv.add_prev\[0\] VSS VSS VCC VCC _0574_ sky130_fd_sc_hd__and2_1
X_4338_ _1964_ _1965_ VSS VSS VCC VCC _1966_ sky130_fd_sc_hd__or2_1
X_4269_ _1895_ _1896_ VSS VSS VCC VCC _1897_ sky130_fd_sc_hd__or2_1
X_3640_ _0807_ _1411_ _1522_ VSS VSS VCC VCC _1523_ sky130_fd_sc_hd__o21ai_1
X_3571_ _1458_ _1457_ net184 net354 VSS VSS VCC VCC _1459_ sky130_fd_sc_hd__a2bb2o_1
X_2522_ _0492_ _0493_ _0495_ VSS VSS VCC VCC _0497_ sky130_fd_sc_hd__a21o_1
X_5310_ clknet_leaf_168_i_clk _0338_ VSS VSS VCC VCC u_muldiv.dividend\[25\]
+ sky130_fd_sc_hd__dfxtp_4
X_2453_ net590 VSS VSS VCC VCC _0428_ sky130_fd_sc_hd__inv_2
X_5241_ clknet_leaf_126_i_clk _0269_ VSS VSS VCC VCC u_muldiv.o_div\[18\]
+ sky130_fd_sc_hd__dfxtp_2
X_5172_ clknet_4_12__leaf_i_clk _0204_ VSS VSS VCC VCC u_muldiv.add_prev\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_4123_ net583 net582 _1816_ net382 VSS VSS VCC VCC _1824_ sky130_fd_sc_hd__o31a_1
X_4054_ net592 _1768_ _1769_ VSS VSS VCC VCC _1770_ sky130_fd_sc_hd__o21ba_1
Xinput2 i_alu_ctrl[1] VSS VSS VCC VCC net2 sky130_fd_sc_hd__buf_8
X_3005_ u_muldiv.dividend\[26\] net419 net364 u_muldiv.o_div\[26\] net442 vssd1 vssd1
+ vccd1 vccd1 _0971_ sky130_fd_sc_hd__a221o_1
X_4956_ _1210_ net400 VSS VSS VCC VCC _0400_ sky130_fd_sc_hd__nor2_1
X_3907_ net501 net101 net723 VSS VSS VCC VCC _1712_ sky130_fd_sc_hd__and3_1
X_4887_ net571 _2422_ net459 net650 VSS VSS VCC VCC _2423_ sky130_fd_sc_hd__o211a_1
X_3838_ net592 net723 _1660_ _1659_ VSS VSS VCC VCC _0057_ sky130_fd_sc_hd__o22a_1
X_3769_ net502 net241 net723 _1612_ VSS VSS VCC VCC _0036_ sky130_fd_sc_hd__o211a_1
X_4810_ net480 _2352_ VSS VSS VCC VCC _2353_ sky130_fd_sc_hd__nor2_1
X_4741_ _2266_ _2289_ VSS VSS VCC VCC _2290_ sky130_fd_sc_hd__nand2_1
X_4672_ net697 net695 _2207_ VSS VSS VCC VCC _2227_ sky130_fd_sc_hd__or3_2
X_3623_ _1119_ net606 _0766_ _1506_ VSS VSS VCC VCC _1507_ sky130_fd_sc_hd__a211o_1
X_3554_ u_bits.i_op2\[9\] net699 net353 VSS VSS VCC VCC _1443_ sky130_fd_sc_hd__a21oi_1
X_2505_ _0477_ _0478_ _0479_ VSS VSS VCC VCC _0480_ sky130_fd_sc_hd__nand3_2
X_3485_ net575 u_pc_sel.i_pc_next\[4\] _1377_ _1378_ VSS VSS VCC VCC net271
+ sky130_fd_sc_hd__a22o_4
X_5224_ clknet_leaf_93_i_clk _0252_ VSS VSS VCC VCC u_muldiv.o_div\[1\] sky130_fd_sc_hd__dfxtp_2
X_5155_ clknet_leaf_68_i_clk _0187_ VSS VSS VCC VCC u_muldiv.add_prev\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4106_ net585 _1810_ net384 VSS VSS VCC VCC _1811_ sky130_fd_sc_hd__o21ai_1
X_5086_ clknet_leaf_60_i_clk _0119_ VSS VSS VCC VCC net290 sky130_fd_sc_hd__dfxtp_4
X_4037_ u_muldiv.divisor\[40\] net483 net335 u_muldiv.divisor\[41\] _1756_ vssd1 vssd1
+ vccd1 vccd1 _0160_ sky130_fd_sc_hd__a221o_1
Xclkbuf_4_1__f_i_clk clknet_2_0_0_i_clk VSS VSS VCC VCC clknet_4_1__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4939_ _1166_ _1169_ net406 VSS VSS VCC VCC _0383_ sky130_fd_sc_hd__and3_1
Xoutput191 net191 VSS VSS VCC VCC o_add[17] sky130_fd_sc_hd__buf_2
Xclkbuf_2_2_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_2_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_3270_ _0499_ _1207_ VSS VSS VCC VCC _1208_ sky130_fd_sc_hd__xnor2_4
X_2985_ net663 net584 net410 _0951_ _0952_ VSS VSS VCC VCC _0953_ sky130_fd_sc_hd__a311oi_2
X_4724_ _1916_ _1918_ _2272_ VSS VSS VCC VCC _2274_ sky130_fd_sc_hd__a21o_1
X_4655_ u_muldiv.dividend\[10\] net324 net375 _2211_ VSS VSS VCC VCC _0323_
+ sky130_fd_sc_hd__a31o_1
Xinput60 i_op1[23] VSS VSS VCC VCC net60 sky130_fd_sc_hd__clkbuf_1
X_3606_ net574 u_pc_sel.i_pc_next\[12\] _1490_ _1491_ VSS VSS VCC VCC net248
+ sky130_fd_sc_hd__a22o_4
Xclkbuf_leaf_6_i_clk clknet_4_1__leaf_i_clk VSS VSS VCC VCC clknet_leaf_6_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput71 i_op1[4] VSS VSS VCC VCC net71 sky130_fd_sc_hd__clkbuf_1
X_4586_ net438 _2142_ _2146_ _2147_ _2148_ VSS VSS VCC VCC _2149_ sky130_fd_sc_hd__a32o_1
Xinput82 i_op2[14] VSS VSS VCC VCC net82 sky130_fd_sc_hd__clkbuf_4
Xinput93 i_op2[24] VSS VSS VCC VCC net93 sky130_fd_sc_hd__clkbuf_1
X_3537_ _1270_ _1271_ _1275_ _1276_ net619 net450 VSS VSS VCC VCC _1427_ sky130_fd_sc_hd__mux4_1
X_3468_ net619 _1271_ VSS VSS VCC VCC _1362_ sky130_fd_sc_hd__or2_1
X_5207_ clknet_leaf_157_i_clk _0239_ VSS VSS VCC VCC u_muldiv.mul\[24\] sky130_fd_sc_hd__dfxtp_1
X_3399_ _0933_ _1295_ net450 VSS VSS VCC VCC _1296_ sky130_fd_sc_hd__mux2_1
X_5138_ clknet_leaf_42_i_clk _0170_ VSS VSS VCC VCC u_muldiv.divisor\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_5069_ clknet_leaf_134_i_clk _0102_ VSS VSS VCC VCC net234 sky130_fd_sc_hd__dfxtp_4
X_2770_ _0744_ _0533_ _0528_ VSS VSS VCC VCC _0745_ sky130_fd_sc_hd__a21oi_4
X_4440_ u_muldiv.quotient_msk\[16\] u_muldiv.o_div\[16\] net470 net436 vssd1 vssd1
+ vccd1 vccd1 _2053_ sky130_fd_sc_hd__o211a_1
X_4371_ net470 net491 net376 VSS VSS VCC VCC _1998_ sky130_fd_sc_hd__o21a_2
X_3322_ _1251_ net561 VSS VSS VCC VCC _1252_ sky130_fd_sc_hd__nand2_1
Xfanout609 net610 VSS VSS VCC VCC net609 sky130_fd_sc_hd__buf_6
X_3253_ _0646_ _1193_ _0660_ VSS VSS VCC VCC _1195_ sky130_fd_sc_hd__a21o_1
X_3184_ _1140_ VSS VSS VCC VCC net207 sky130_fd_sc_hd__clkinv_4
X_2968_ _0935_ VSS VSS VCC VCC _0936_ sky130_fd_sc_hd__inv_2
X_4707_ u_muldiv.dividend\[14\] _2239_ u_muldiv.dividend\[15\] VSS VSS VCC VCC
+ _2259_ sky130_fd_sc_hd__o21ai_1
X_2899_ u_muldiv.mul\[56\] net363 net357 u_muldiv.mul\[24\] VSS VSS VCC VCC
+ _0870_ sky130_fd_sc_hd__a22oi_1
Xclkbuf_leaf_154_i_clk clknet_4_9__leaf_i_clk VSS VSS VCC VCC clknet_leaf_154_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4638_ net704 net702 _2172_ net373 net699 VSS VSS VCC VCC _2196_ sky130_fd_sc_hd__o311a_1
X_4569_ _2131_ net374 net712 VSS VSS VCC VCC _2133_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_107_i_clk clknet_4_9__leaf_i_clk VSS VSS VCC VCC clknet_leaf_107_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3940_ net220 net124 net386 VSS VSS VCC VCC _0103_ sky130_fd_sc_hd__mux2_1
X_3871_ net586 u_bits.i_op2\[21\] net546 VSS VSS VCC VCC _1685_ sky130_fd_sc_hd__mux2_1
X_2822_ net612 _0795_ net606 VSS VSS VCC VCC _0796_ sky130_fd_sc_hd__o21ai_1
X_2753_ _0706_ _0726_ VSS VSS VCC VCC _0728_ sky130_fd_sc_hd__nor2_1
X_2684_ net428 _0652_ _0653_ _0657_ VSS VSS VCC VCC _0659_ sky130_fd_sc_hd__a31o_2
X_4423_ _2035_ u_muldiv.o_div\[13\] net492 net385 VSS VSS VCC VCC _2039_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_86_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_86_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4354_ u_muldiv.divisor\[55\] u_muldiv.divisor\[54\] u_muldiv.divisor\[53\] u_muldiv.divisor\[52\]
+ VSS VSS VCC VCC _1982_ sky130_fd_sc_hd__or4_1
Xfanout406 net407 VSS VSS VCC VCC net406 sky130_fd_sc_hd__buf_4
Xfanout417 net418 VSS VSS VCC VCC net417 sky130_fd_sc_hd__buf_4
Xfanout428 net430 VSS VSS VCC VCC net428 sky130_fd_sc_hd__buf_6
X_3305_ _0832_ _1225_ _1230_ _1234_ VSS VSS VCC VCC _1235_ sky130_fd_sc_hd__nand4_1
Xfanout439 _0451_ VSS VSS VCC VCC net439 sky130_fd_sc_hd__buf_12
X_4285_ u_muldiv.divisor\[16\] u_muldiv.dividend\[16\] VSS VSS VCC VCC _1913_
+ sky130_fd_sc_hd__and2b_1
X_3236_ _1181_ VSS VSS VCC VCC net214 sky130_fd_sc_hd__inv_2
X_3167_ _0422_ _1123_ _1124_ net206 net355 VSS VSS VCC VCC _1125_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_24_i_clk clknet_4_6__leaf_i_clk VSS VSS VCC VCC clknet_leaf_24_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3098_ _1037_ _1038_ _1059_ VSS VSS VCC VCC _1060_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_39_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_39_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4070_ _1781_ _1782_ VSS VSS VCC VCC _1783_ sky130_fd_sc_hd__nor2_1
X_3021_ net661 u_bits.i_op2\[26\] net410 _0986_ VSS VSS VCC VCC _0987_ sky130_fd_sc_hd__a31o_1
X_4972_ clknet_leaf_43_i_clk _0005_ VSS VSS VCC VCC u_bits.i_op1\[2\] sky130_fd_sc_hd__dfxtp_4
X_3923_ u_pc_sel.i_pc_next\[14\] net113 net391 VSS VSS VCC VCC _0089_ sky130_fd_sc_hd__mux2_1
X_3854_ net589 net727 _1672_ _1671_ VSS VSS VCC VCC _0061_ sky130_fd_sc_hd__o22a_1
X_2805_ _0778_ VSS VSS VCC VCC _0779_ sky130_fd_sc_hd__inv_2
X_3785_ net505 net545 net725 net626 VSS VSS VCC VCC _1621_ sky130_fd_sc_hd__and4bb_1
X_2736_ net703 u_muldiv.add_prev\[8\] net540 VSS VSS VCC VCC _0711_ sky130_fd_sc_hd__mux2_1
X_2667_ _0640_ _0641_ net432 VSS VSS VCC VCC _0642_ sky130_fd_sc_hd__nand3_1
X_4406_ net318 _2025_ u_muldiv.o_div\[9\] VSS VSS VCC VCC _2026_ sky130_fd_sc_hd__a21oi_1
X_2598_ _0419_ net537 _0572_ VSS VSS VCC VCC _0573_ sky130_fd_sc_hd__o21ai_1
X_4337_ u_muldiv.dividend\[28\] u_muldiv.divisor\[28\] VSS VSS VCC VCC _1965_
+ sky130_fd_sc_hd__and2b_1
X_4268_ _0445_ u_muldiv.divisor\[12\] VSS VSS VCC VCC _1896_ sky130_fd_sc_hd__and2_1
X_3219_ _1167_ _1168_ VSS VSS VCC VCC net210 sky130_fd_sc_hd__nand2_8
X_4199_ u_muldiv.mul\[29\] u_muldiv.mul\[28\] net405 VSS VSS VCC VCC _0243_
+ sky130_fd_sc_hd__mux2_1
X_3570_ net352 _1452_ _1455_ _1456_ net521 VSS VSS VCC VCC _1458_ sky130_fd_sc_hd__a41o_1
X_2521_ _0492_ _0493_ _0495_ VSS VSS VCC VCC _0496_ sky130_fd_sc_hd__a21oi_1
X_5240_ clknet_leaf_126_i_clk _0268_ VSS VSS VCC VCC u_muldiv.o_div\[17\]
+ sky130_fd_sc_hd__dfxtp_2
X_2452_ net596 VSS VSS VCC VCC _0427_ sky130_fd_sc_hd__inv_2
X_5171_ clknet_leaf_61_i_clk _0203_ VSS VSS VCC VCC u_muldiv.add_prev\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_4122_ net583 net582 _1816_ VSS VSS VCC VCC _1823_ sky130_fd_sc_hd__or3_1
X_4053_ net592 _1768_ net486 net468 VSS VSS VCC VCC _1769_ sky130_fd_sc_hd__a211o_1
Xinput3 i_alu_ctrl[2] VSS VSS VCC VCC net3 sky130_fd_sc_hd__clkbuf_1
X_3004_ _0970_ VSS VSS VCC VCC net201 sky130_fd_sc_hd__inv_6
X_4955_ net555 net195 _0432_ VSS VSS VCC VCC _0399_ sky130_fd_sc_hd__and3b_1
X_3906_ net580 net728 _1711_ _1710_ VSS VSS VCC VCC _0074_ sky130_fd_sc_hd__o22a_1
X_4886_ net656 net654 net652 _2388_ VSS VSS VCC VCC _2422_ sky130_fd_sc_hd__nor4_1
X_3837_ net501 net81 net720 VSS VSS VCC VCC _1660_ sky130_fd_sc_hd__a21o_1
X_3768_ net176 net501 VSS VSS VCC VCC _1612_ sky130_fd_sc_hd__nand2b_1
X_2719_ _0692_ _0691_ _0689_ VSS VSS VCC VCC _0694_ sky130_fd_sc_hd__nand3b_2
X_3699_ net409 _1574_ _1577_ _1572_ VSS VSS VCC VCC _1578_ sky130_fd_sc_hd__o211a_1
X_5369_ clknet_leaf_152_i_clk _0396_ VSS VSS VCC VCC u_muldiv.mul\[48\] sky130_fd_sc_hd__dfxtp_1
X_4740_ net684 net682 VSS VSS VCC VCC _2289_ sky130_fd_sc_hd__nor2_1
X_4671_ _1892_ _1895_ _1896_ net470 VSS VSS VCC VCC _2226_ sky130_fd_sc_hd__o31a_1
X_3622_ _0772_ _0857_ _1395_ _0806_ VSS VSS VCC VCC _1506_ sky130_fd_sc_hd__a2bb2o_1
X_3553_ net596 net699 net351 _1441_ VSS VSS VCC VCC _1442_ sky130_fd_sc_hd__o211ai_1
X_2504_ net674 u_muldiv.add_prev\[21\] net531 VSS VSS VCC VCC _0479_ sky130_fd_sc_hd__mux2_1
X_3484_ net32 net730 net574 VSS VSS VCC VCC _1378_ sky130_fd_sc_hd__o21ba_1
X_5223_ clknet_leaf_100_i_clk net500 VSS VSS VCC VCC u_muldiv.on_wait sky130_fd_sc_hd__dfxtp_4
X_5154_ clknet_leaf_67_i_clk _0186_ VSS VSS VCC VCC u_muldiv.add_prev\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4105_ net586 _1806_ net379 VSS VSS VCC VCC _1810_ sky130_fd_sc_hd__o21ai_1
X_5085_ clknet_leaf_144_i_clk _0118_ VSS VSS VCC VCC net279 sky130_fd_sc_hd__dfxtp_4
X_4036_ net596 _1754_ _1755_ VSS VSS VCC VCC _1756_ sky130_fd_sc_hd__a21oi_1
X_4938_ _1162_ _1163_ net401 VSS VSS VCC VCC _0382_ sky130_fd_sc_hd__a21oi_2
X_4869_ _2406_ _2405_ _2401_ _2403_ VSS VSS VCC VCC _2407_ sky130_fd_sc_hd__o22a_1
Xoutput192 net192 VSS VSS VCC VCC o_add[18] sky130_fd_sc_hd__buf_2
X_2984_ net601 _0934_ net327 VSS VSS VCC VCC _0952_ sky130_fd_sc_hd__o21a_1
X_4723_ _2272_ _1916_ VSS VSS VCC VCC _2273_ sky130_fd_sc_hd__nand2_1
X_4654_ net494 _2205_ _2210_ net318 _2202_ VSS VSS VCC VCC _2211_ sky130_fd_sc_hd__o311a_1
X_3605_ net9 net730 net574 VSS VSS VCC VCC _1491_ sky130_fd_sc_hd__o21ba_1
Xinput50 i_op1[14] VSS VSS VCC VCC net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 i_op1[24] VSS VSS VCC VCC net61 sky130_fd_sc_hd__clkbuf_1
Xinput72 i_op1[5] VSS VSS VCC VCC net72 sky130_fd_sc_hd__clkbuf_1
X_4585_ _0444_ _2136_ net497 VSS VSS VCC VCC _2148_ sky130_fd_sc_hd__o21a_1
Xinput83 i_op2[15] VSS VSS VCC VCC net83 sky130_fd_sc_hd__buf_2
Xinput94 i_op2[25] VSS VSS VCC VCC net94 sky130_fd_sc_hd__buf_4
X_3536_ _0894_ net601 VSS VSS VCC VCC _1426_ sky130_fd_sc_hd__nand2b_1
X_3467_ net346 _1273_ _1275_ _0905_ _1360_ VSS VSS VCC VCC _1361_ sky130_fd_sc_hd__o221a_1
X_5206_ clknet_leaf_157_i_clk _0238_ VSS VSS VCC VCC u_muldiv.mul\[23\] sky130_fd_sc_hd__dfxtp_1
X_3398_ _1293_ _1294_ net619 VSS VSS VCC VCC _1295_ sky130_fd_sc_hd__mux2_1
X_5137_ clknet_leaf_42_i_clk _0169_ VSS VSS VCC VCC u_muldiv.divisor\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_5068_ clknet_leaf_82_i_clk _0101_ VSS VSS VCC VCC net233 sky130_fd_sc_hd__dfxtp_1
X_4019_ net603 net600 _1279_ net382 VSS VSS VCC VCC _1742_ sky130_fd_sc_hd__o31a_1
X_4370_ u_muldiv.o_div\[1\] _1997_ net321 VSS VSS VCC VCC _0252_ sky130_fd_sc_hd__mux2_1
X_3321_ _1250_ _1247_ _1249_ VSS VSS VCC VCC _1251_ sky130_fd_sc_hd__o21ai_1
X_3252_ _0649_ _1192_ _0660_ _0646_ VSS VSS VCC VCC _1194_ sky130_fd_sc_hd__o211ai_4
X_3183_ _1138_ _1139_ VSS VSS VCC VCC _1140_ sky130_fd_sc_hd__nand2_2
X_2967_ net628 _0847_ VSS VSS VCC VCC _0935_ sky130_fd_sc_hd__or2_1
X_4706_ u_muldiv.dividend\[15\] u_muldiv.dividend\[14\] u_muldiv.dividend\[13\] _2222_
+ VSS VSS VCC VCC _2258_ sky130_fd_sc_hd__or4_2
X_2898_ u_muldiv.dividend\[24\] net419 net364 u_muldiv.o_div\[24\] vssd1 vssd1 vccd1
+ vccd1 _0869_ sky130_fd_sc_hd__a22oi_1
X_4637_ net704 net702 _2172_ net372 VSS VSS VCC VCC _2195_ sky130_fd_sc_hd__o31a_1
X_4568_ net461 net718 net716 net713 net374 VSS VSS VCC VCC _2132_ sky130_fd_sc_hd__o311a_1
X_3519_ _1340_ _1343_ net456 VSS VSS VCC VCC _1410_ sky130_fd_sc_hd__mux2_1
X_4499_ _2095_ net477 u_muldiv.o_div\[29\] net383 VSS VSS VCC VCC _2099_ sky130_fd_sc_hd__a31o_1
X_3870_ u_bits.i_op2\[21\] net725 _1684_ _1683_ VSS VSS VCC VCC _0065_ sky130_fd_sc_hd__o22a_1
X_2821_ _0788_ _0790_ _0793_ _0791_ net629 net620 VSS VSS VCC VCC _0795_ sky130_fd_sc_hd__mux4_2
X_2752_ _0726_ VSS VSS VCC VCC _0727_ sky130_fd_sc_hd__inv_2
X_2683_ _0655_ _0656_ _0657_ VSS VSS VCC VCC _0658_ sky130_fd_sc_hd__o21ai_4
X_4422_ u_muldiv.o_div\[12\] _2038_ net318 VSS VSS VCC VCC _0263_ sky130_fd_sc_hd__mux2_1
X_4353_ u_muldiv.divisor\[35\] u_muldiv.divisor\[34\] u_muldiv.divisor\[33\] u_muldiv.divisor\[32\]
+ VSS VSS VCC VCC _1981_ sky130_fd_sc_hd__or4_1
Xfanout407 net408 VSS VSS VCC VCC net407 sky130_fd_sc_hd__buf_6
X_3304_ _1030_ _1036_ _1233_ _1210_ _1201_ VSS VSS VCC VCC _1234_ sky130_fd_sc_hd__o2111a_1
Xfanout418 _0757_ VSS VSS VCC VCC net418 sky130_fd_sc_hd__buf_12
Xfanout429 net430 VSS VSS VCC VCC net429 sky130_fd_sc_hd__clkbuf_4
X_4284_ _1910_ _1911_ VSS VSS VCC VCC _1912_ sky130_fd_sc_hd__nand2_1
X_3235_ _1179_ _1180_ VSS VSS VCC VCC _1181_ sky130_fd_sc_hd__nand2_2
X_3166_ net653 net580 net440 _0781_ VSS VSS VCC VCC _1124_ sky130_fd_sc_hd__a211o_1
X_3097_ _1058_ _1057_ net203 net355 net527 VSS VSS VCC VCC _1059_ sky130_fd_sc_hd__a221o_1
X_3999_ _1725_ _1726_ net330 VSS VSS VCC VCC _1727_ sky130_fd_sc_hd__a21oi_1
X_3020_ _0979_ _0901_ net345 _0983_ VSS VSS VCC VCC _0986_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_153_i_clk clknet_4_8__leaf_i_clk VSS VSS VCC VCC clknet_leaf_153_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4971_ clknet_leaf_48_i_clk _0004_ VSS VSS VCC VCC u_bits.i_op1\[1\] sky130_fd_sc_hd__dfxtp_4
X_3922_ u_pc_sel.i_pc_next\[13\] net112 net392 VSS VSS VCC VCC _0088_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_168_i_clk clknet_4_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_168_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3853_ net512 net85 net721 VSS VSS VCC VCC _1672_ sky130_fd_sc_hd__a21o_1
X_2804_ _0772_ _0777_ net615 VSS VSS VCC VCC _0778_ sky130_fd_sc_hd__mux2_1
X_3784_ net505 net77 net725 VSS VSS VCC VCC _1620_ sky130_fd_sc_hd__and3_1
X_2735_ net518 net526 _0707_ _0708_ VSS VSS VCC VCC _0710_ sky130_fd_sc_hd__o211ai_2
X_2666_ net448 net593 VSS VSS VCC VCC _0641_ sky130_fd_sc_hd__nand2_1
X_4405_ _2020_ u_muldiv.quotient_msk\[9\] net435 VSS VSS VCC VCC _2025_ sky130_fd_sc_hd__mux2_1
X_5385_ clknet_leaf_90_i_clk _0412_ VSS VSS VCC VCC u_bits.i_op1\[0\] sky130_fd_sc_hd__dfxtp_2
X_2597_ net648 net555 _0571_ net425 VSS VSS VCC VCC _0572_ sky130_fd_sc_hd__o211ai_2
X_4336_ u_muldiv.divisor\[28\] u_muldiv.dividend\[28\] VSS VSS VCC VCC _1964_
+ sky130_fd_sc_hd__and2b_1
X_4267_ u_muldiv.divisor\[12\] _0445_ VSS VSS VCC VCC _1895_ sky130_fd_sc_hd__nor2_2
X_3218_ _0591_ _0600_ _0601_ _1166_ VSS VSS VCC VCC _1168_ sky130_fd_sc_hd__nand4_4
X_4198_ u_muldiv.mul\[28\] u_muldiv.mul\[27\] net405 VSS VSS VCC VCC _0242_
+ sky130_fd_sc_hd__mux2_1
X_3149_ _1106_ _1107_ VSS VSS VCC VCC _1108_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_70_i_clk clknet_4_13__leaf_i_clk VSS VSS VCC VCC clknet_leaf_70_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_85_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_85_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2520_ net446 net678 _0494_ VSS VSS VCC VCC _0495_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_23_i_clk clknet_4_6__leaf_i_clk VSS VSS VCC VCC clknet_leaf_23_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2451_ net598 VSS VSS VCC VCC _0426_ sky130_fd_sc_hd__inv_4
X_5170_ clknet_leaf_72_i_clk _0202_ VSS VSS VCC VCC u_muldiv.add_prev\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_4121_ u_muldiv.divisor\[58\] net482 net337 u_muldiv.divisor\[59\] _1822_ vssd1 vssd1
+ vccd1 vccd1 _0178_ sky130_fd_sc_hd__a221o_1
X_4052_ net594 net593 _1760_ net381 VSS VSS VCC VCC _1768_ sky130_fd_sc_hd__o31a_1
Xinput4 i_alu_ctrl[3] VSS VSS VCC VCC net4 sky130_fd_sc_hd__clkbuf_1
X_3003_ _0967_ _0969_ VSS VSS VCC VCC _0970_ sky130_fd_sc_hd__xnor2_4
X_4954_ _1208_ net402 VSS VSS VCC VCC _0398_ sky130_fd_sc_hd__nor2_2
X_3905_ net513 net100 net721 VSS VSS VCC VCC _1711_ sky130_fd_sc_hd__a21o_1
X_4885_ _1973_ _2420_ VSS VSS VCC VCC _2421_ sky130_fd_sc_hd__nand2_1
X_3836_ net503 _1658_ VSS VSS VCC VCC _1659_ sky130_fd_sc_hd__and2b_1
X_3767_ net501 net277 net723 _1611_ VSS VSS VCC VCC _0035_ sky130_fd_sc_hd__o211a_1
X_2718_ _0688_ _0690_ _0692_ VSS VSS VCC VCC _0693_ sky130_fd_sc_hd__o21ai_4
X_3698_ net587 net678 net411 _1576_ VSS VSS VCC VCC _1577_ sky130_fd_sc_hd__a31oi_4
X_2649_ net448 net707 _0622_ VSS VSS VCC VCC _0624_ sky130_fd_sc_hd__a21oi_1
X_5368_ clknet_leaf_76_i_clk _0395_ VSS VSS VCC VCC u_muldiv.mul\[47\] sky130_fd_sc_hd__dfxtp_2
X_4319_ u_muldiv.divisor\[25\] u_muldiv.dividend\[25\] VSS VSS VCC VCC _1947_
+ sky130_fd_sc_hd__xnor2_2
X_5299_ clknet_leaf_142_i_clk _0327_ VSS VSS VCC VCC u_muldiv.dividend\[14\]
+ sky130_fd_sc_hd__dfxtp_4
Xfanout590 u_bits.i_op2\[16\] VSS VSS VCC VCC net590 sky130_fd_sc_hd__clkbuf_8
X_4670_ _1897_ _1892_ VSS VSS VCC VCC _2225_ sky130_fd_sc_hd__nor2_1
X_3621_ _1505_ u_pc_sel.i_pc_next\[13\] net576 VSS VSS VCC VCC net249 sky130_fd_sc_hd__mux2_8
X_3552_ _0427_ net569 net700 VSS VSS VCC VCC _1441_ sky130_fd_sc_hd__or3b_1
X_2503_ net517 net523 _0476_ VSS VSS VCC VCC _0478_ sky130_fd_sc_hd__o21ai_1
X_3483_ net443 _1373_ _1376_ net733 VSS VSS VCC VCC _1377_ sky130_fd_sc_hd__a211o_2
X_5222_ clknet_leaf_45_i_clk _0251_ VSS VSS VCC VCC op_cnt\[5\] sky130_fd_sc_hd__dfxtp_1
X_5153_ clknet_leaf_67_i_clk _0185_ VSS VSS VCC VCC u_muldiv.add_prev\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4104_ u_muldiv.divisor\[54\] net484 net335 u_muldiv.divisor\[55\] _1809_ vssd1 vssd1
+ vccd1 vccd1 _0174_ sky130_fd_sc_hd__a221o_1
X_5084_ clknet_leaf_21_i_clk _0117_ VSS VSS VCC VCC net278 sky130_fd_sc_hd__dfxtp_4
X_4035_ net596 _1754_ net384 VSS VSS VCC VCC _1755_ sky130_fd_sc_hd__o21ai_1
X_4937_ _1165_ net402 VSS VSS VCC VCC _0381_ sky130_fd_sc_hd__nor2_1
X_4868_ _2404_ net369 net654 net330 VSS VSS VCC VCC _2406_ sky130_fd_sc_hd__a31o_1
X_3819_ net595 net597 net548 VSS VSS VCC VCC _1646_ sky130_fd_sc_hd__mux2_1
X_4799_ u_muldiv.dividend\[22\] _2322_ u_muldiv.dividend\[23\] VSS VSS VCC VCC
+ _2343_ sky130_fd_sc_hd__o21ai_1
Xoutput193 net193 VSS VSS VCC VCC o_add[19] sky130_fd_sc_hd__buf_2
X_2983_ net662 net584 _0950_ net348 VSS VSS VCC VCC _0951_ sky130_fd_sc_hd__o211a_1
X_4722_ _1908_ _1915_ _1913_ VSS VSS VCC VCC _2272_ sky130_fd_sc_hd__a21oi_1
X_4653_ net697 _2208_ _2209_ VSS VSS VCC VCC _2210_ sky130_fd_sc_hd__o21ba_1
Xinput40 i_funct3[0] VSS VSS VCC VCC net40 sky130_fd_sc_hd__clkbuf_4
X_3604_ net527 _1486_ _1489_ net730 VSS VSS VCC VCC _1490_ sky130_fd_sc_hd__o211ai_4
Xinput51 i_op1[15] VSS VSS VCC VCC net51 sky130_fd_sc_hd__clkbuf_1
X_4584_ u_muldiv.dividend\[3\] u_muldiv.dividend\[4\] _2126_ VSS VSS VCC VCC
+ _2147_ sky130_fd_sc_hd__or3_1
Xinput62 i_op1[25] VSS VSS VCC VCC net62 sky130_fd_sc_hd__buf_2
Xinput73 i_op1[6] VSS VSS VCC VCC net73 sky130_fd_sc_hd__clkbuf_1
Xinput84 i_op2[16] VSS VSS VCC VCC net84 sky130_fd_sc_hd__buf_6
Xinput95 i_op2[26] VSS VSS VCC VCC net95 sky130_fd_sc_hd__buf_2
X_3535_ u_bits.i_op2\[8\] net701 _1424_ net350 VSS VSS VCC VCC _1425_ sky130_fd_sc_hd__o211ai_1
X_3466_ net611 _1359_ VSS VSS VCC VCC _1360_ sky130_fd_sc_hd__nand2_1
X_5205_ clknet_leaf_159_i_clk _0237_ VSS VSS VCC VCC u_muldiv.mul\[22\] sky130_fd_sc_hd__dfxtp_1
X_3397_ net670 net665 net672 net668 net625 net458 VSS VSS VCC VCC _1294_ sky130_fd_sc_hd__mux4_2
X_5136_ clknet_4_5__leaf_i_clk _0168_ VSS VSS VCC VCC u_muldiv.divisor\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_5067_ clknet_leaf_81_i_clk _0100_ VSS VSS VCC VCC net232 sky130_fd_sc_hd__dfxtp_2
X_4018_ _0806_ _0840_ net456 _0425_ VSS VSS VCC VCC _1741_ sky130_fd_sc_hd__nand4_4
X_3320_ u_adder.i_cmp_inverse _1135_ VSS VSS VCC VCC _1250_ sky130_fd_sc_hd__nand2b_1
X_3251_ _0736_ _1191_ _0650_ VSS VSS VCC VCC _1193_ sky130_fd_sc_hd__o21ai_4
X_3182_ _1108_ _1101_ _1106_ _1137_ VSS VSS VCC VCC _1139_ sky130_fd_sc_hd__o211ai_4
X_2966_ net612 _0933_ net347 VSS VSS VCC VCC _0934_ sky130_fd_sc_hd__o21a_1
X_4705_ net469 _2253_ _2256_ net488 VSS VSS VCC VCC _2257_ sky130_fd_sc_hd__a211oi_1
X_2897_ net731 net21 _0868_ VSS VSS VCC VCC net260 sky130_fd_sc_hd__o21a_2
X_4636_ u_muldiv.dividend\[7\] u_muldiv.dividend\[9\] u_muldiv.dividend\[8\] _2161_
+ VSS VSS VCC VCC _2194_ sky130_fd_sc_hd__nor4_4
X_4567_ net460 net718 net716 VSS VSS VCC VCC _2131_ sky130_fd_sc_hd__or3_2
X_3518_ net578 u_pc_sel.i_pc_next\[6\] _1408_ _1409_ VSS VSS VCC VCC net273
+ sky130_fd_sc_hd__a22o_2
X_4498_ u_muldiv.o_div\[28\] _2098_ net315 VSS VSS VCC VCC _0279_ sky130_fd_sc_hd__mux2_1
X_3449_ _0905_ _1343_ net609 VSS VSS VCC VCC _1344_ sky130_fd_sc_hd__o21ba_1
X_5119_ clknet_leaf_6_i_clk _0151_ VSS VSS VCC VCC u_muldiv.divisor\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_2820_ _0793_ _0791_ net629 VSS VSS VCC VCC _0794_ sky130_fd_sc_hd__mux2_1
X_2751_ _0713_ _0714_ _0724_ _0725_ VSS VSS VCC VCC _0726_ sky130_fd_sc_hd__nand4_4
X_2682_ net692 u_muldiv.add_prev\[13\] net542 VSS VSS VCC VCC _0657_ sky130_fd_sc_hd__mux2_1
X_4421_ _2036_ net493 _2035_ _2037_ VSS VSS VCC VCC _2038_ sky130_fd_sc_hd__a31o_1
X_4352_ u_muldiv.divisor\[43\] u_muldiv.divisor\[42\] u_muldiv.divisor\[41\] u_muldiv.divisor\[40\]
+ VSS VSS VCC VCC _1980_ sky130_fd_sc_hd__or4_1
Xfanout408 _1255_ VSS VSS VCC VCC net408 sky130_fd_sc_hd__buf_6
X_3303_ _1030_ _1036_ u_adder.i_cmp_inverse VSS VSS VCC VCC _1233_ sky130_fd_sc_hd__a21boi_1
X_4283_ u_muldiv.dividend\[19\] u_muldiv.divisor\[19\] VSS VSS VCC VCC _1911_
+ sky130_fd_sc_hd__nand2b_1
Xfanout419 net422 VSS VSS VCC VCC net419 sky130_fd_sc_hd__buf_4
X_3234_ _0712_ _1178_ _0725_ _0724_ VSS VSS VCC VCC _1180_ sky130_fd_sc_hd__o211ai_2
X_3165_ net410 _1117_ _1120_ _1122_ VSS VSS VCC VCC _1123_ sky130_fd_sc_hd__or4_1
X_3096_ net410 _1053_ net522 VSS VSS VCC VCC _1058_ sky130_fd_sc_hd__a21oi_1
X_3998_ net640 net378 net626 VSS VSS VCC VCC _1726_ sky130_fd_sc_hd__a21bo_1
X_2949_ net22 net729 VSS VSS VCC VCC _0919_ sky130_fd_sc_hd__nor2_1
X_4619_ _2176_ _2178_ net322 VSS VSS VCC VCC _2179_ sky130_fd_sc_hd__a21oi_1
X_4970_ net461 net45 net398 VSS VSS VCC VCC _0412_ sky130_fd_sc_hd__mux2_1
X_3921_ u_pc_sel.i_pc_next\[12\] net111 net396 VSS VSS VCC VCC _0087_ sky130_fd_sc_hd__mux2_1
X_3852_ net512 _1670_ VSS VSS VCC VCC _1671_ sky130_fd_sc_hd__and2b_1
X_2803_ net622 _0776_ _0773_ VSS VSS VCC VCC _0777_ sky130_fd_sc_hd__o21a_1
X_3783_ net515 u_pc_sel.i_inst_branch net728 _1619_ VSS VSS VCC VCC _0043_
+ sky130_fd_sc_hd__o211a_1
X_2734_ _0707_ _0708_ net428 VSS VSS VCC VCC _0709_ sky130_fd_sc_hd__a21o_1
X_2665_ net647 net552 _0639_ net424 VSS VSS VCC VCC _0640_ sky130_fd_sc_hd__o211ai_2
X_4404_ _2020_ u_muldiv.o_div\[9\] net492 net385 VSS VSS VCC VCC _2024_ sky130_fd_sc_hd__a31o_1
X_2596_ net537 net460 VSS VSS VCC VCC _0571_ sky130_fd_sc_hd__and2_1
X_5384_ clknet_leaf_23_i_clk _0411_ VSS VSS VCC VCC u_muldiv.mul\[63\] sky130_fd_sc_hd__dfxtp_1
X_4335_ u_muldiv.dividend\[29\] u_muldiv.divisor\[29\] VSS VSS VCC VCC _1963_
+ sky130_fd_sc_hd__nand2b_1
X_4266_ u_muldiv.divisor\[13\] u_muldiv.dividend\[13\] VSS VSS VCC VCC _1894_
+ sky130_fd_sc_hd__xor2_1
X_3217_ _0600_ _0601_ _1166_ _0591_ VSS VSS VCC VCC _1167_ sky130_fd_sc_hd__a22o_2
X_4197_ u_muldiv.mul\[27\] u_muldiv.mul\[26\] net405 VSS VSS VCC VCC _0241_
+ sky130_fd_sc_hd__mux2_1
X_3148_ _1104_ _1103_ VSS VSS VCC VCC _1107_ sky130_fd_sc_hd__or2_1
X_3079_ net615 _1039_ net347 VSS VSS VCC VCC _1041_ sky130_fd_sc_hd__o21ai_1
X_2450_ net600 VSS VSS VCC VCC _0425_ sky130_fd_sc_hd__inv_6
X_4120_ _1820_ _1821_ net383 VSS VSS VCC VCC _1822_ sky130_fd_sc_hd__and3_1
X_4051_ u_muldiv.divisor\[43\] net484 net335 u_muldiv.divisor\[44\] _1767_ vssd1 vssd1
+ vccd1 vccd1 _0163_ sky130_fd_sc_hd__a221o_1
Xinput5 i_alu_ctrl[4] VSS VSS VCC VCC net5 sky130_fd_sc_hd__clkbuf_1
X_3002_ _0888_ _0927_ _0877_ _0968_ VSS VSS VCC VCC _0969_ sky130_fd_sc_hd__a31oi_4
X_4953_ net555 net192 _0432_ VSS VSS VCC VCC _0397_ sky130_fd_sc_hd__and3b_1
X_3904_ net515 _1709_ VSS VSS VCC VCC _1710_ sky130_fd_sc_hd__and2b_1
X_4884_ _1974_ _1984_ u_muldiv.divisor\[30\] _0447_ VSS VSS VCC VCC _2420_
+ sky130_fd_sc_hd__o2bb2a_1
X_3835_ u_bits.i_op2\[14\] net593 net545 VSS VSS VCC VCC _1658_ sky130_fd_sc_hd__mux2_1
X_3766_ net181 net501 VSS VSS VCC VCC _1611_ sky130_fd_sc_hd__nand2b_1
X_2717_ net698 u_muldiv.add_prev\[10\] net540 VSS VSS VCC VCC _0692_ sky130_fd_sc_hd__mux2_1
X_3697_ net587 net678 _1575_ net349 VSS VSS VCC VCC _1576_ sky130_fd_sc_hd__o211a_1
X_2648_ net448 net707 VSS VSS VCC VCC _0623_ sky130_fd_sc_hd__and2_1
X_5367_ clknet_4_12__leaf_i_clk _0394_ VSS VSS VCC VCC u_muldiv.mul\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_2579_ _0548_ _0550_ net428 VSS VSS VCC VCC _0554_ sky130_fd_sc_hd__a21oi_2
X_4318_ u_muldiv.divisor\[24\] u_muldiv.dividend\[24\] VSS VSS VCC VCC _1946_
+ sky130_fd_sc_hd__xnor2_2
X_5298_ clknet_4_8__leaf_i_clk _0326_ VSS VSS VCC VCC u_muldiv.dividend\[13\]
+ sky130_fd_sc_hd__dfxtp_4
X_4249_ u_muldiv.dividend\[8\] u_muldiv.divisor\[8\] VSS VSS VCC VCC _1877_
+ sky130_fd_sc_hd__nand2b_1
Xclkbuf_leaf_152_i_clk clknet_4_9__leaf_i_clk VSS VSS VCC VCC clknet_leaf_152_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_167_i_clk clknet_4_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_167_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout580 u_bits.i_op2\[30\] VSS VSS VCC VCC net580 sky130_fd_sc_hd__buf_6
Xfanout591 u_bits.i_op2\[15\] VSS VSS VCC VCC net591 sky130_fd_sc_hd__clkbuf_8
X_3620_ _1504_ net10 net734 VSS VSS VCC VCC _1505_ sky130_fd_sc_hd__mux2_2
X_3551_ _1438_ _1439_ _0910_ _0941_ VSS VSS VCC VCC _1440_ sky130_fd_sc_hd__o2bb2a_2
X_2502_ net531 _0431_ net432 _0475_ VSS VSS VCC VCC _0477_ sky130_fd_sc_hd__o211ai_2
X_3482_ net556 u_muldiv.mul\[4\] net415 net529 _1375_ VSS VSS VCC VCC _1376_
+ sky130_fd_sc_hd__o311a_1
X_5221_ clknet_leaf_49_i_clk _0250_ VSS VSS VCC VCC op_cnt\[4\] sky130_fd_sc_hd__dfxtp_1
X_5152_ clknet_leaf_103_i_clk _0184_ VSS VSS VCC VCC u_muldiv.add_prev\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4103_ _1807_ _1808_ VSS VSS VCC VCC _1809_ sky130_fd_sc_hd__nor2_1
X_5083_ clknet_leaf_59_i_clk _0116_ VSS VSS VCC VCC u_mux.i_add_override sky130_fd_sc_hd__dfxtp_2
X_4034_ net598 net597 _1745_ net379 VSS VSS VCC VCC _1754_ sky130_fd_sc_hd__o31a_1
X_4936_ net402 _1213_ VSS VSS VCC VCC _0380_ sky130_fd_sc_hd__nor2_1
X_4867_ _2404_ net370 net654 VSS VSS VCC VCC _2405_ sky130_fd_sc_hd__a21oi_1
X_3818_ net597 net728 _1645_ _1644_ VSS VSS VCC VCC _0052_ sky130_fd_sc_hd__o22a_1
X_4798_ u_muldiv.dividend\[23\] u_muldiv.dividend\[22\] _2322_ VSS VSS VCC VCC
+ _2342_ sky130_fd_sc_hd__or3_2
X_3749_ net687 net51 net396 VSS VSS VCC VCC _0018_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_84_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_84_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xoutput183 net183 VSS VSS VCC VCC o_add[0] sky130_fd_sc_hd__buf_2
Xoutput194 net194 VSS VSS VCC VCC o_add[1] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_22_i_clk clknet_4_6__leaf_i_clk VSS VSS VCC VCC clknet_leaf_22_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_37_i_clk clknet_4_4__leaf_i_clk VSS VSS VCC VCC clknet_leaf_37_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2982_ net560 net584 net662 VSS VSS VCC VCC _0950_ sky130_fd_sc_hd__nand3b_1
X_4721_ u_muldiv.dividend\[16\] net326 net377 _2271_ VSS VSS VCC VCC _0329_
+ sky130_fd_sc_hd__a31o_1
X_4652_ _2207_ net372 net697 net472 VSS VSS VCC VCC _2209_ sky130_fd_sc_hd__a31o_1
X_3603_ net557 u_muldiv.mul\[12\] net413 net528 _1488_ VSS VSS VCC VCC _1489_
+ sky130_fd_sc_hd__o311ai_4
Xinput30 i_csr_data[31] VSS VSS VCC VCC net30 sky130_fd_sc_hd__buf_4
Xinput41 i_funct3[1] VSS VSS VCC VCC net41 sky130_fd_sc_hd__buf_4
Xinput52 i_op1[16] VSS VSS VCC VCC net52 sky130_fd_sc_hd__clkbuf_1
X_4583_ net711 _2144_ _2145_ VSS VSS VCC VCC _2146_ sky130_fd_sc_hd__o21ai_1
Xinput63 i_op1[26] VSS VSS VCC VCC net63 sky130_fd_sc_hd__clkbuf_1
Xinput74 i_op1[7] VSS VSS VCC VCC net74 sky130_fd_sc_hd__clkbuf_1
Xinput85 i_op2[17] VSS VSS VCC VCC net85 sky130_fd_sc_hd__clkbuf_4
X_3534_ net567 net701 net597 VSS VSS VCC VCC _1424_ sky130_fd_sc_hd__nand3b_1
Xinput96 i_op2[27] VSS VSS VCC VCC net96 sky130_fd_sc_hd__buf_2
X_3465_ net619 _1276_ _1358_ VSS VSS VCC VCC _1359_ sky130_fd_sc_hd__o21ai_1
X_5204_ clknet_leaf_160_i_clk _0236_ VSS VSS VCC VCC u_muldiv.mul\[21\] sky130_fd_sc_hd__dfxtp_1
X_3396_ net682 net679 net677 net675 net642 net631 VSS VSS VCC VCC _1293_ sky130_fd_sc_hd__mux4_2
X_5135_ clknet_leaf_39_i_clk _0167_ VSS VSS VCC VCC u_muldiv.divisor\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_5066_ clknet_leaf_72_i_clk _0099_ VSS VSS VCC VCC net231 sky130_fd_sc_hd__dfxtp_1
X_4017_ u_muldiv.divisor\[36\] net482 net337 u_muldiv.divisor\[37\] _1740_ vssd1 vssd1
+ vccd1 vccd1 _0156_ sky130_fd_sc_hd__a221o_1
X_4919_ u_muldiv.divisor\[26\] net475 net332 u_muldiv.divisor\[27\] vssd1 vssd1 vccd1
+ vccd1 _0371_ sky130_fd_sc_hd__a22o_1
X_3250_ _0638_ _0728_ _0736_ VSS VSS VCC VCC _1192_ sky130_fd_sc_hd__a21oi_2
X_3181_ _1105_ _1109_ _1137_ VSS VSS VCC VCC _1138_ sky130_fd_sc_hd__o21bai_2
X_2965_ _0932_ _0931_ net619 VSS VSS VCC VCC _0933_ sky130_fd_sc_hd__mux2_1
X_4704_ net686 _2254_ _2255_ VSS VSS VCC VCC _2256_ sky130_fd_sc_hd__o21a_1
X_2896_ net577 _0867_ VSS VSS VCC VCC _0868_ sky130_fd_sc_hd__nor2_1
X_4635_ u_muldiv.dividend\[7\] u_muldiv.dividend\[8\] _2161_ u_muldiv.dividend\[9\]
+ VSS VSS VCC VCC _2193_ sky130_fd_sc_hd__o31a_1
X_4566_ _1852_ _1854_ _1862_ VSS VSS VCC VCC _2130_ sky130_fd_sc_hd__or3_1
X_3517_ net34 net731 net577 VSS VSS VCC VCC _1409_ sky130_fd_sc_hd__o21ba_1
X_4497_ _2095_ _2096_ net477 _2097_ VSS VSS VCC VCC _2098_ sky130_fd_sc_hd__a31o_1
X_3448_ net705 net703 net700 net698 net646 net634 VSS VSS VCC VCC _1343_ sky130_fd_sc_hd__mux4_1
X_3379_ _1273_ _1274_ _1276_ _1275_ net454 net614 VSS VSS VCC VCC _1277_ sky130_fd_sc_hd__mux4_1
X_5118_ clknet_leaf_58_i_clk mul_op2_signed_next VSS VSS VCC VCC u_muldiv.i_op2_signed
+ sky130_fd_sc_hd__dfxtp_1
X_5049_ clknet_leaf_129_i_clk _0082_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_2750_ _0720_ _0721_ _0718_ _0719_ VSS VSS VCC VCC _0725_ sky130_fd_sc_hd__o211ai_4
X_2681_ _0652_ _0653_ net428 VSS VSS VCC VCC _0656_ sky130_fd_sc_hd__a21oi_4
X_4420_ u_muldiv.quotient_msk\[12\] u_muldiv.o_div\[12\] net471 net435 vssd1 vssd1
+ vccd1 vccd1 _2037_ sky130_fd_sc_hd__o211a_1
X_4351_ u_muldiv.divisor\[39\] u_muldiv.divisor\[38\] u_muldiv.divisor\[37\] u_muldiv.divisor\[36\]
+ VSS VSS VCC VCC _1979_ sky130_fd_sc_hd__or4_1
X_3302_ _1222_ _1231_ u_adder.i_cmp_inverse VSS VSS VCC VCC _1232_ sky130_fd_sc_hd__o21bai_1
Xfanout409 _0815_ VSS VSS VCC VCC net409 sky130_fd_sc_hd__clkbuf_8
X_4282_ u_muldiv.divisor\[19\] u_muldiv.dividend\[19\] VSS VSS VCC VCC _1910_
+ sky130_fd_sc_hd__nand2b_1
X_3233_ _0724_ _0725_ _0638_ _0714_ _0712_ VSS VSS VCC VCC _1179_ sky130_fd_sc_hd__a221o_1
X_3164_ net653 net580 _1121_ net348 VSS VSS VCC VCC _1122_ sky130_fd_sc_hd__o211a_1
X_3095_ net410 _1042_ _1055_ _1056_ VSS VSS VCC VCC _1057_ sky130_fd_sc_hd__or4_1
X_3997_ net458 net626 net570 net579 VSS VSS VCC VCC _1725_ sky130_fd_sc_hd__or4b_1
X_2948_ net527 _0869_ _0870_ _0917_ VSS VSS VCC VCC _0918_ sky130_fd_sc_hd__a31o_1
X_2879_ net616 _0850_ net608 VSS VSS VCC VCC _0851_ sky130_fd_sc_hd__o21ai_1
X_4618_ u_muldiv.dividend\[7\] _2161_ _2177_ VSS VSS VCC VCC _2178_ sky130_fd_sc_hd__a21o_1
X_4549_ net461 net717 net374 VSS VSS VCC VCC _2115_ sky130_fd_sc_hd__and3_1
X_3920_ u_pc_sel.i_pc_next\[11\] net110 net388 VSS VSS VCC VCC _0086_ sky130_fd_sc_hd__mux2_1
X_3851_ net588 net590 net548 VSS VSS VCC VCC _1670_ sky130_fd_sc_hd__mux2_1
X_2802_ net632 _0775_ _0774_ VSS VSS VCC VCC _0776_ sky130_fd_sc_hd__o21a_1
X_3782_ net43 net515 VSS VSS VCC VCC _1619_ sky130_fd_sc_hd__nand2b_1
X_2733_ net449 u_bits.i_op2\[8\] VSS VSS VCC VCC _0708_ sky130_fd_sc_hd__nand2_1
X_2664_ net542 net694 VSS VSS VCC VCC _0639_ sky130_fd_sc_hd__and2_1
X_4403_ u_muldiv.o_div\[8\] _2023_ net320 VSS VSS VCC VCC _0259_ sky130_fd_sc_hd__mux2_1
X_5383_ clknet_leaf_19_i_clk _0410_ VSS VSS VCC VCC u_muldiv.mul\[62\] sky130_fd_sc_hd__dfxtp_1
X_2595_ net447 net648 VSS VSS VCC VCC _0570_ sky130_fd_sc_hd__nand2_1
X_4334_ u_muldiv.divisor\[29\] u_muldiv.dividend\[29\] VSS VSS VCC VCC _1962_
+ sky130_fd_sc_hd__nand2b_1
X_4265_ _1884_ _1889_ _1891_ VSS VSS VCC VCC _1893_ sky130_fd_sc_hd__o21bai_1
X_3216_ _0582_ _0583_ _0593_ VSS VSS VCC VCC _1166_ sky130_fd_sc_hd__a21o_2
X_4196_ u_muldiv.mul\[26\] u_muldiv.mul\[25\] net405 VSS VSS VCC VCC _0240_
+ sky130_fd_sc_hd__mux2_1
X_3147_ _1105_ VSS VSS VCC VCC _1106_ sky130_fd_sc_hd__clkinv_2
X_3078_ net611 _1039_ net347 VSS VSS VCC VCC _1040_ sky130_fd_sc_hd__o21a_1
Xclkbuf_4_4__f_i_clk clknet_2_1_0_i_clk VSS VSS VCC VCC clknet_4_4__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4050_ _1765_ _1766_ VSS VSS VCC VCC _1767_ sky130_fd_sc_hd__nor2_1
X_3001_ _0875_ _0926_ _0925_ VSS VSS VCC VCC _0968_ sky130_fd_sc_hd__o21ai_2
Xinput6 i_csr_data[0] VSS VSS VCC VCC net6 sky130_fd_sc_hd__clkbuf_2
X_4952_ net400 _1221_ VSS VSS VCC VCC _0396_ sky130_fd_sc_hd__nor2_2
X_3903_ net579 net581 net549 VSS VSS VCC VCC _1709_ sky130_fd_sc_hd__mux2_1
X_4883_ _1843_ _1972_ _1974_ _1984_ VSS VSS VCC VCC _2419_ sky130_fd_sc_hd__o211ai_1
X_3834_ net593 net727 _1657_ _1656_ VSS VSS VCC VCC _0056_ sky130_fd_sc_hd__o22a_1
X_3765_ u_bits.i_op1\[31\] net69 net387 VSS VSS VCC VCC _0034_ sky130_fd_sc_hd__mux2_1
X_2716_ net518 net525 _0686_ _0687_ VSS VSS VCC VCC _0691_ sky130_fd_sc_hd__o211ai_1
X_3696_ net561 net678 net587 VSS VSS VCC VCC _1575_ sky130_fd_sc_hd__nand3b_1
Xoutput310 net310 VSS VSS VCC VCC o_wdata[9] sky130_fd_sc_hd__buf_2
X_2647_ net540 u_muldiv.add_prev\[6\] VSS VSS VCC VCC _0622_ sky130_fd_sc_hd__and2_1
X_5366_ clknet_leaf_75_i_clk _0393_ VSS VSS VCC VCC u_muldiv.mul\[45\] sky130_fd_sc_hd__dfxtp_2
X_2578_ net518 net525 _0551_ VSS VSS VCC VCC _0553_ sky130_fd_sc_hd__o21ai_2
X_4317_ u_muldiv.divisor\[24\] u_muldiv.dividend\[24\] VSS VSS VCC VCC _1945_
+ sky130_fd_sc_hd__nand2b_1
X_5297_ clknet_4_9__leaf_i_clk _0325_ VSS VSS VCC VCC u_muldiv.dividend\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_4248_ u_muldiv.divisor\[8\] u_muldiv.dividend\[8\] VSS VSS VCC VCC _1876_
+ sky130_fd_sc_hd__nand2b_1
X_4179_ u_muldiv.mul\[9\] u_muldiv.mul\[8\] net403 VSS VSS VCC VCC _0223_
+ sky130_fd_sc_hd__mux2_1
Xfanout570 net571 VSS VSS VCC VCC net570 sky130_fd_sc_hd__buf_6
Xfanout581 u_bits.i_op2\[29\] VSS VSS VCC VCC net581 sky130_fd_sc_hd__buf_6
Xfanout592 u_bits.i_op2\[13\] VSS VSS VCC VCC net592 sky130_fd_sc_hd__buf_8
X_3550_ _0857_ _1295_ _1299_ _0807_ _0765_ VSS VSS VCC VCC _1439_ sky130_fd_sc_hd__o221a_1
X_2501_ net531 _0431_ _0475_ VSS VSS VCC VCC _0476_ sky130_fd_sc_hd__o21ai_1
X_3481_ u_muldiv.o_div\[4\] net366 net358 _1374_ VSS VSS VCC VCC _1375_ sky130_fd_sc_hd__a211o_1
X_5220_ clknet_leaf_45_i_clk _0249_ VSS VSS VCC VCC op_cnt\[3\] sky130_fd_sc_hd__dfxtp_1
X_5151_ clknet_leaf_9_i_clk _0183_ VSS VSS VCC VCC u_muldiv.quotient_msk\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_4102_ _1806_ net380 net586 net329 VSS VSS VCC VCC _1808_ sky130_fd_sc_hd__a31o_1
X_5082_ clknet_leaf_8_i_clk _0115_ VSS VSS VCC VCC u_bits.i_sra sky130_fd_sc_hd__dfxtp_4
X_4033_ net599 net598 net597 _1741_ VSS VSS VCC VCC _1753_ sky130_fd_sc_hd__nor4_1
Xclkbuf_leaf_3_i_clk clknet_4_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_3_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4935_ _0576_ _1211_ net406 VSS VSS VCC VCC _0379_ sky130_fd_sc_hd__and3_1
X_4866_ net658 net656 _2338_ _2379_ VSS VSS VCC VCC _2404_ sky130_fd_sc_hd__or4b_1
X_3817_ net512 net107 net721 VSS VSS VCC VCC _1645_ sky130_fd_sc_hd__a21o_1
X_4797_ net480 _2339_ _2340_ _1720_ VSS VSS VCC VCC _2341_ sky130_fd_sc_hd__o31ai_1
X_3748_ net688 net50 net395 VSS VSS VCC VCC _0017_ sky130_fd_sc_hd__mux2_1
X_3679_ net601 _1320_ net327 VSS VSS VCC VCC _1559_ sky130_fd_sc_hd__o21a_1
X_5349_ clknet_leaf_23_i_clk _0003_ VSS VSS VCC VCC u_muldiv.add_prev\[31\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput184 net184 VSS VSS VCC VCC o_add[10] sky130_fd_sc_hd__buf_2
Xoutput195 net195 VSS VSS VCC VCC o_add[20] sky130_fd_sc_hd__buf_2
X_2981_ _0945_ net611 _0948_ VSS VSS VCC VCC _0949_ sky130_fd_sc_hd__a21bo_1
X_4720_ _2265_ _2270_ net319 _2263_ VSS VSS VCC VCC _2271_ sky130_fd_sc_hd__o211a_1
X_4651_ net701 net699 _2184_ net372 VSS VSS VCC VCC _2208_ sky130_fd_sc_hd__o31a_1
Xinput20 i_csr_data[22] VSS VSS VCC VCC net20 sky130_fd_sc_hd__buf_4
X_3602_ u_muldiv.o_div\[12\] net366 net358 _1487_ VSS VSS VCC VCC _1488_ sky130_fd_sc_hd__a211o_1
Xinput31 i_csr_data[3] VSS VSS VCC VCC net31 sky130_fd_sc_hd__buf_4
X_4582_ _2144_ net711 net474 VSS VSS VCC VCC _2145_ sky130_fd_sc_hd__a21oi_1
Xinput42 i_funct3[2] VSS VSS VCC VCC net42 sky130_fd_sc_hd__buf_6
Xinput53 i_op1[17] VSS VSS VCC VCC net53 sky130_fd_sc_hd__clkbuf_1
Xinput64 i_op1[27] VSS VSS VCC VCC net64 sky130_fd_sc_hd__clkbuf_1
Xinput75 i_op1[8] VSS VSS VCC VCC net75 sky130_fd_sc_hd__clkbuf_1
X_3533_ net243 u_pc_sel.i_pc_next\[7\] _1422_ _1423_ VSS VSS VCC VCC net274
+ sky130_fd_sc_hd__a22o_4
Xinput86 i_op2[18] VSS VSS VCC VCC net86 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput97 i_op2[28] VSS VSS VCC VCC net97 sky130_fd_sc_hd__clkbuf_1
X_3464_ net453 _1270_ VSS VSS VCC VCC _1358_ sky130_fd_sc_hd__or2_1
X_5203_ clknet_leaf_151_i_clk _0235_ VSS VSS VCC VCC u_muldiv.mul\[20\] sky130_fd_sc_hd__dfxtp_1
X_3395_ net731 _1291_ _1292_ VSS VSS VCC VCC net245 sky130_fd_sc_hd__a21oi_2
X_5134_ clknet_leaf_39_i_clk _0166_ VSS VSS VCC VCC u_muldiv.divisor\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_5065_ clknet_leaf_0_i_clk _0098_ VSS VSS VCC VCC net230 sky130_fd_sc_hd__dfxtp_1
X_4016_ _0425_ _1738_ _1739_ VSS VSS VCC VCC _1740_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_151_i_clk clknet_4_9__leaf_i_clk VSS VSS VCC VCC clknet_leaf_151_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4918_ u_muldiv.divisor\[25\] net476 net332 u_muldiv.divisor\[26\] vssd1 vssd1 vccd1
+ vccd1 _0370_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_166_i_clk clknet_4_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_166_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4849_ net658 _2338_ _2379_ VSS VSS VCC VCC _2388_ sky130_fd_sc_hd__or3b_2
Xclkbuf_leaf_104_i_clk clknet_4_12__leaf_i_clk VSS VSS VCC VCC clknet_leaf_104_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_119_i_clk clknet_4_11__leaf_i_clk VSS VSS VCC VCC clknet_leaf_119_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3180_ _1135_ _1136_ VSS VSS VCC VCC _1137_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_83_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_83_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2964_ net663 net660 net658 net656 net637 net625 VSS VSS VCC VCC _0932_ sky130_fd_sc_hd__mux4_2
X_4703_ _2254_ net686 net469 VSS VSS VCC VCC _2255_ sky130_fd_sc_hd__a21oi_1
X_2895_ _0834_ _0866_ net735 VSS VSS VCC VCC _0867_ sky130_fd_sc_hd__a21oi_4
X_4634_ _2190_ _2191_ net459 net494 VSS VSS VCC VCC _2192_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_98_i_clk clknet_4_12__leaf_i_clk VSS VSS VCC VCC clknet_leaf_98_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4565_ _1852_ _1854_ _1862_ VSS VSS VCC VCC _2129_ sky130_fd_sc_hd__o21ai_1
X_3516_ net444 _1404_ _1407_ net734 VSS VSS VCC VCC _1408_ sky130_fd_sc_hd__a211o_1
X_4496_ u_muldiv.quotient_msk\[28\] u_muldiv.o_div\[28\] net465 net433 vssd1 vssd1
+ vccd1 vccd1 _2097_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_21_i_clk clknet_4_3__leaf_i_clk VSS VSS VCC VCC clknet_leaf_21_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3447_ net712 net711 net708 net707 net646 net635 VSS VSS VCC VCC _1342_ sky130_fd_sc_hd__mux4_1
X_3378_ net693 net690 net688 net686 net643 net630 VSS VSS VCC VCC _1276_ sky130_fd_sc_hd__mux4_2
X_5117_ clknet_leaf_24_i_clk _0150_ VSS VSS VCC VCC u_adder.i_cmp_inverse
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_36_i_clk clknet_4_4__leaf_i_clk VSS VSS VCC VCC clknet_leaf_36_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5048_ clknet_leaf_78_i_clk _0081_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_2680_ _0463_ _0651_ _0654_ VSS VSS VCC VCC _0655_ sky130_fd_sc_hd__a21oi_2
X_4350_ u_muldiv.divisor\[59\] u_muldiv.divisor\[58\] u_muldiv.divisor\[57\] u_muldiv.divisor\[56\]
+ VSS VSS VCC VCC _1978_ sky130_fd_sc_hd__or4_2
X_3301_ _1223_ _1225_ _1230_ _1140_ VSS VSS VCC VCC _1231_ sky130_fd_sc_hd__nand4_1
X_4281_ u_muldiv.divisor\[18\] u_muldiv.dividend\[18\] VSS VSS VCC VCC _1909_
+ sky130_fd_sc_hd__xor2_1
X_3232_ _0636_ _0637_ _0715_ VSS VSS VCC VCC _1178_ sky130_fd_sc_hd__a21oi_1
X_3163_ net561 net580 net653 VSS VSS VCC VCC _1121_ sky130_fd_sc_hd__nand3b_1
X_3094_ _1047_ _0814_ net601 _1052_ VSS VSS VCC VCC _1056_ sky130_fd_sc_hd__a31o_1
X_3996_ net570 net579 VSS VSS VCC VCC _1724_ sky130_fd_sc_hd__and2b_1
X_2947_ _0422_ _0916_ net199 net355 net527 VSS VSS VCC VCC _0917_ sky130_fd_sc_hd__a221oi_4
X_2878_ net457 _0848_ _0849_ VSS VSS VCC VCC _0850_ sky130_fd_sc_hd__o21ai_2
X_4617_ u_muldiv.dividend\[7\] _2161_ net494 VSS VSS VCC VCC _2177_ sky130_fd_sc_hd__o21ai_1
X_4548_ net573 net650 VSS VSS VCC VCC _2114_ sky130_fd_sc_hd__nand2b_4
X_4479_ _2081_ _2082_ net481 _2083_ VSS VSS VCC VCC _2084_ sky130_fd_sc_hd__a31o_1
X_3850_ net590 net726 _1669_ _1668_ VSS VSS VCC VCC _0060_ sky130_fd_sc_hd__o22a_1
X_2801_ net652 net650 net639 VSS VSS VCC VCC _0775_ sky130_fd_sc_hd__mux2_1
X_3781_ net515 u_pc_sel.i_inst_jal_jalr net728 _1618_ VSS VSS VCC VCC _0042_
+ sky130_fd_sc_hd__o211a_1
X_2732_ net648 net554 net703 net540 net426 VSS VSS VCC VCC _0707_ sky130_fd_sc_hd__o2111ai_2
X_2663_ _0636_ _0637_ VSS VSS VCC VCC _0638_ sky130_fd_sc_hd__nand2_2
X_4402_ _2020_ _2021_ net493 _2022_ VSS VSS VCC VCC _2023_ sky130_fd_sc_hd__a31o_1
X_2594_ _0565_ _0566_ _0567_ VSS VSS VCC VCC _0569_ sky130_fd_sc_hd__nand3_1
X_5382_ clknet_leaf_23_i_clk _0409_ VSS VSS VCC VCC u_muldiv.mul\[61\] sky130_fd_sc_hd__dfxtp_1
X_4333_ u_muldiv.divisor\[29\] u_muldiv.dividend\[29\] VSS VSS VCC VCC _1961_
+ sky130_fd_sc_hd__and2b_1
X_4264_ _1884_ _1889_ _1891_ VSS VSS VCC VCC _1892_ sky130_fd_sc_hd__o21ba_1
X_3215_ _1165_ VSS VSS VCC VCC net205 sky130_fd_sc_hd__inv_4
X_4195_ u_muldiv.mul\[25\] u_muldiv.mul\[24\] net405 VSS VSS VCC VCC _0239_
+ sky130_fd_sc_hd__mux2_1
X_3146_ _1103_ _1104_ VSS VSS VCC VCC _1105_ sky130_fd_sc_hd__and2_1
X_3077_ net619 _0892_ _0773_ VSS VSS VCC VCC _1039_ sky130_fd_sc_hd__o21a_1
X_3979_ u_wr_mux.i_reg_data2\[23\] net159 net387 VSS VSS VCC VCC _0141_ sky130_fd_sc_hd__mux2_1
Xfanout730 net732 VSS VSS VCC VCC net730 sky130_fd_sc_hd__buf_6
X_3000_ _0964_ _0965_ VSS VSS VCC VCC _0967_ sky130_fd_sc_hd__nand2_2
Xinput7 i_csr_data[10] VSS VSS VCC VCC net7 sky130_fd_sc_hd__clkbuf_4
X_4951_ _1205_ _1218_ net406 VSS VSS VCC VCC _0395_ sky130_fd_sc_hd__and3_1
X_3902_ net581 net727 _1708_ _1707_ VSS VSS VCC VCC _0073_ sky130_fd_sc_hd__o22a_1
X_4882_ u_muldiv.dividend\[30\] net315 _2418_ VSS VSS VCC VCC _0343_ sky130_fd_sc_hd__o21a_1
X_3833_ net510 net80 net721 VSS VSS VCC VCC _1657_ sky130_fd_sc_hd__a21o_1
X_3764_ net653 net68 net396 VSS VSS VCC VCC _0033_ sky130_fd_sc_hd__mux2_1
X_2715_ net519 net525 _0686_ _0687_ VSS VSS VCC VCC _0690_ sky130_fd_sc_hd__o211a_1
X_3695_ _1013_ _0806_ _1009_ _0856_ _1573_ VSS VSS VCC VCC _1574_ sky130_fd_sc_hd__a221o_1
Xoutput300 net300 VSS VSS VCC VCC o_wdata[29] sky130_fd_sc_hd__buf_2
X_2646_ net518 net525 _0616_ _0617_ VSS VSS VCC VCC _0621_ sky130_fd_sc_hd__o211ai_1
Xoutput311 net311 VSS VSS VCC VCC o_wsel[0] sky130_fd_sc_hd__buf_2
X_5365_ clknet_leaf_77_i_clk _0392_ VSS VSS VCC VCC u_muldiv.mul\[44\] sky130_fd_sc_hd__dfxtp_2
X_2577_ net457 net537 _0460_ _0549_ net432 VSS VSS VCC VCC _0552_ sky130_fd_sc_hd__o221ai_4
X_4316_ _1941_ _1925_ _1943_ VSS VSS VCC VCC _1944_ sky130_fd_sc_hd__o21bai_4
X_5296_ clknet_leaf_155_i_clk _0324_ VSS VSS VCC VCC u_muldiv.dividend\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_4247_ _1873_ _1866_ _1846_ _1870_ VSS VSS VCC VCC _1875_ sky130_fd_sc_hd__o211a_1
X_4178_ net736 u_muldiv.mul\[7\] net403 VSS VSS VCC VCC _0222_ sky130_fd_sc_hd__mux2_1
X_3129_ _0905_ _0946_ net346 _1088_ net345 VSS VSS VCC VCC _1089_ sky130_fd_sc_hd__o221ai_1
Xfanout560 net561 VSS VSS VCC VCC net560 sky130_fd_sc_hd__buf_4
Xfanout571 net215 VSS VSS VCC VCC net571 sky130_fd_sc_hd__buf_6
Xfanout582 u_bits.i_op2\[27\] VSS VSS VCC VCC net582 sky130_fd_sc_hd__buf_4
Xfanout593 u_bits.i_op2\[12\] VSS VSS VCC VCC net593 sky130_fd_sc_hd__buf_8
X_2500_ net646 net551 net532 net674 net423 VSS VSS VCC VCC _0475_ sky130_fd_sc_hd__o2111ai_2
X_3480_ net568 net558 u_muldiv.dividend\[4\] u_muldiv.mul\[36\] net362 vssd1 vssd1
+ vccd1 vccd1 _1374_ sky130_fd_sc_hd__a32o_1
X_5150_ clknet_leaf_10_i_clk _0182_ VSS VSS VCC VCC u_muldiv.divisor\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_4101_ _1806_ net380 net586 VSS VSS VCC VCC _1807_ sky130_fd_sc_hd__a21oi_1
X_5081_ clknet_leaf_73_i_clk _0114_ VSS VSS VCC VCC alu_ctrl\[2\] sky130_fd_sc_hd__dfxtp_2
X_4032_ u_muldiv.divisor\[39\] net482 net335 u_muldiv.divisor\[40\] _1752_ vssd1 vssd1
+ vccd1 vccd1 _0159_ sky130_fd_sc_hd__a221o_1
X_4934_ u_muldiv.dividend\[0\] _2435_ _1989_ VSS VSS VCC VCC _0378_ sky130_fd_sc_hd__mux2_1
X_4865_ _2402_ net476 VSS VSS VCC VCC _2403_ sky130_fd_sc_hd__nand2_1
X_3816_ net513 _1643_ VSS VSS VCC VCC _1644_ sky130_fd_sc_hd__and2b_1
X_4796_ _2338_ net369 net667 VSS VSS VCC VCC _2340_ sky130_fd_sc_hd__a21oi_1
X_3747_ net692 net49 net395 VSS VSS VCC VCC _0016_ sky130_fd_sc_hd__mux2_1
X_3678_ u_muldiv.mul\[50\] net361 net360 u_muldiv.mul\[18\] _1557_ vssd1 vssd1 vccd1
+ vccd1 _1558_ sky130_fd_sc_hd__a221o_1
X_2629_ _0591_ _0592_ _0600_ _0601_ VSS VSS VCC VCC _0604_ sky130_fd_sc_hd__nand4_1
X_5348_ clknet_leaf_22_i_clk _0376_ VSS VSS VCC VCC u_muldiv.outsign sky130_fd_sc_hd__dfxtp_2
Xoutput185 net185 VSS VSS VCC VCC o_add[11] sky130_fd_sc_hd__buf_2
Xoutput196 net196 VSS VSS VCC VCC o_add[21] sky130_fd_sc_hd__buf_2
X_5279_ clknet_4_0__leaf_i_clk _0307_ VSS VSS VCC VCC u_muldiv.quotient_msk\[24\]
+ sky130_fd_sc_hd__dfxtp_2
Xfanout390 net391 VSS VSS VCC VCC net390 sky130_fd_sc_hd__clkbuf_4
X_2980_ net346 _0946_ _0947_ _0905_ net345 VSS VSS VCC VCC _0948_ sky130_fd_sc_hd__o221a_1
X_4650_ net704 net701 net699 _2172_ VSS VSS VCC VCC _2207_ sky130_fd_sc_hd__or4_1
X_3601_ net567 net557 u_muldiv.dividend\[12\] u_muldiv.mul\[44\] net362 vssd1 vssd1
+ vccd1 vccd1 _1487_ sky130_fd_sc_hd__a32o_1
Xinput10 i_csr_data[13] VSS VSS VCC VCC net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 i_csr_data[23] VSS VSS VCC VCC net21 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 i_csr_data[4] VSS VSS VCC VCC net32 sky130_fd_sc_hd__clkbuf_4
X_4581_ net713 _2131_ net374 VSS VSS VCC VCC _2144_ sky130_fd_sc_hd__o21ai_1
Xinput43 i_inst_branch VSS VSS VCC VCC net43 sky130_fd_sc_hd__buf_6
Xinput54 i_op1[18] VSS VSS VCC VCC net54 sky130_fd_sc_hd__clkbuf_1
Xinput65 i_op1[28] VSS VSS VCC VCC net65 sky130_fd_sc_hd__clkbuf_1
X_3532_ net35 net731 net577 VSS VSS VCC VCC _1423_ sky130_fd_sc_hd__o21ba_1
Xinput76 i_op1[9] VSS VSS VCC VCC net76 sky130_fd_sc_hd__clkbuf_1
Xinput87 i_op2[19] VSS VSS VCC VCC net87 sky130_fd_sc_hd__buf_4
Xinput98 i_op2[29] VSS VSS VCC VCC net98 sky130_fd_sc_hd__clkbuf_1
X_3463_ _1357_ u_pc_sel.i_pc_next\[3\] net577 VSS VSS VCC VCC net270 sky130_fd_sc_hd__mux2_2
X_5202_ clknet_leaf_151_i_clk _0234_ VSS VSS VCC VCC u_muldiv.mul\[19\] sky130_fd_sc_hd__dfxtp_1
X_3394_ net6 net732 net577 VSS VSS VCC VCC _1292_ sky130_fd_sc_hd__o21bai_2
X_5133_ clknet_leaf_39_i_clk _0165_ VSS VSS VCC VCC u_muldiv.divisor\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_5064_ clknet_leaf_134_i_clk _0097_ VSS VSS VCC VCC net229 sky130_fd_sc_hd__dfxtp_4
X_4015_ _1737_ net379 net600 net329 VSS VSS VCC VCC _1739_ sky130_fd_sc_hd__a31o_1
X_4917_ u_muldiv.divisor\[24\] net476 net333 u_muldiv.divisor\[25\] vssd1 vssd1 vccd1
+ vccd1 _0369_ sky130_fd_sc_hd__a22o_1
X_4848_ _0448_ net323 _2387_ VSS VSS VCC VCC _0340_ sky130_fd_sc_hd__a21oi_1
X_4779_ u_muldiv.dividend\[21\] _2324_ net317 VSS VSS VCC VCC _0334_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_2_i_clk clknet_4_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_2_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2963_ _0839_ _0774_ net632 _0835_ VSS VSS VCC VCC _0931_ sky130_fd_sc_hd__o22a_1
X_4702_ net690 net688 _2234_ net372 VSS VSS VCC VCC _2254_ sky130_fd_sc_hd__o31ai_1
X_2894_ net355 net198 _0865_ _0422_ net544 VSS VSS VCC VCC _0866_ sky130_fd_sc_hd__a221o_1
X_4633_ _1875_ _1878_ _1880_ _1876_ _1844_ VSS VSS VCC VCC _2191_ sky130_fd_sc_hd__o2111ai_1
X_4564_ net463 _2128_ net320 VSS VSS VCC VCC _0315_ sky130_fd_sc_hd__mux2_1
X_3515_ net559 u_muldiv.mul\[6\] net413 net529 _1406_ VSS VSS VCC VCC _1407_
+ sky130_fd_sc_hd__o311a_1
X_4495_ _2094_ u_muldiv.o_div\[28\] VSS VSS VCC VCC _2096_ sky130_fd_sc_hd__nand2_1
X_3446_ _1339_ _1340_ net456 VSS VSS VCC VCC _1341_ sky130_fd_sc_hd__mux2_1
X_3377_ net701 net699 net697 net695 net643 net630 VSS VSS VCC VCC _1275_ sky130_fd_sc_hd__mux4_2
X_5116_ clknet_leaf_83_i_clk _0149_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[31\]
+ sky130_fd_sc_hd__dfxtp_2
X_5047_ clknet_leaf_173_i_clk _0080_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_3300_ net192 net195 _1228_ _1229_ VSS VSS VCC VCC _1230_ sky130_fd_sc_hd__nor4_2
X_4280_ _1906_ _1901_ _1907_ VSS VSS VCC VCC _1908_ sky130_fd_sc_hd__o21bai_4
X_3231_ _1177_ VSS VSS VCC VCC net211 sky130_fd_sc_hd__inv_4
X_3162_ net602 _1118_ net328 VSS VSS VCC VCC _1120_ sky130_fd_sc_hd__o21a_1
X_3093_ net656 u_bits.i_op2\[28\] net348 _1054_ VSS VSS VCC VCC _1055_ sky130_fd_sc_hd__o211a_1
X_3995_ net466 u_muldiv.divisor\[32\] net434 _1723_ VSS VSS VCC VCC _0151_
+ sky130_fd_sc_hd__a31o_1
X_2946_ net665 net585 net410 _0915_ VSS VSS VCC VCC _0916_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_103_i_clk clknet_4_12__leaf_i_clk VSS VSS VCC VCC clknet_leaf_103_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2877_ net623 _0845_ VSS VSS VCC VCC _0849_ sky130_fd_sc_hd__or2_1
X_4616_ _2170_ _2169_ net435 _2175_ VSS VSS VCC VCC _2176_ sky130_fd_sc_hd__o211ai_1
X_4547_ net571 net650 VSS VSS VCC VCC _2113_ sky130_fd_sc_hd__and2b_4
Xclkbuf_leaf_118_i_clk clknet_4_11__leaf_i_clk VSS VSS VCC VCC clknet_leaf_118_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4478_ u_muldiv.quotient_msk\[24\] u_muldiv.o_div\[24\] net467 net434 vssd1 vssd1
+ vccd1 vccd1 _2083_ sky130_fd_sc_hd__o211a_1
X_3429_ net620 net613 _0794_ VSS VSS VCC VCC _1325_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_82_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_82_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_97_i_clk clknet_4_14__leaf_i_clk VSS VSS VCC VCC clknet_leaf_97_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2800_ _0768_ net632 VSS VSS VCC VCC _0774_ sky130_fd_sc_hd__nand2_1
X_3780_ net44 net505 VSS VSS VCC VCC _1618_ sky130_fd_sc_hd__nand2b_1
X_2731_ _0703_ _0700_ _0694_ _0693_ _0702_ VSS VSS VCC VCC _0706_ sky130_fd_sc_hd__o2111ai_4
Xclkbuf_leaf_35_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_35_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2662_ _0628_ _0634_ _0627_ VSS VSS VCC VCC _0637_ sky130_fd_sc_hd__a21boi_4
X_4401_ u_muldiv.quotient_msk\[8\] u_muldiv.o_div\[8\] net471 net435 vssd1 vssd1 vccd1
+ vccd1 _2022_ sky130_fd_sc_hd__o211a_1
X_5381_ clknet_leaf_18_i_clk _0408_ VSS VSS VCC VCC u_muldiv.mul\[60\] sky130_fd_sc_hd__dfxtp_1
X_2593_ _0565_ _0566_ _0567_ VSS VSS VCC VCC _0568_ sky130_fd_sc_hd__a21o_2
X_4332_ _1944_ _1955_ _1959_ VSS VSS VCC VCC _1960_ sky130_fd_sc_hd__a21boi_4
X_4263_ _0416_ u_muldiv.dividend\[11\] _1890_ VSS VSS VCC VCC _1891_ sky130_fd_sc_hd__a21bo_1
X_3214_ _0579_ _1164_ VSS VSS VCC VCC _1165_ sky130_fd_sc_hd__nand2_2
X_4194_ u_muldiv.mul\[24\] u_muldiv.mul\[23\] net405 VSS VSS VCC VCC _0238_
+ sky130_fd_sc_hd__mux2_1
X_3145_ net652 u_muldiv.add_prev\[30\] net532 VSS VSS VCC VCC _1104_ sky130_fd_sc_hd__mux2_1
X_3076_ u_muldiv.mul\[60\] net363 net357 u_muldiv.mul\[28\] VSS VSS VCC VCC
+ _1038_ sky130_fd_sc_hd__a22o_1
X_3978_ u_wr_mux.i_reg_data2\[22\] net158 net390 VSS VSS VCC VCC _0140_ sky130_fd_sc_hd__mux2_1
X_2929_ _0798_ _0790_ _0788_ _0793_ net620 net629 VSS VSS VCC VCC _0899_ sky130_fd_sc_hd__mux4_2
Xfanout720 net722 VSS VSS VCC VCC net720 sky130_fd_sc_hd__buf_4
Xfanout731 net732 VSS VSS VCC VCC net731 sky130_fd_sc_hd__buf_8
Xinput8 i_csr_data[11] VSS VSS VCC VCC net8 sky130_fd_sc_hd__clkbuf_2
X_4950_ _1201_ net402 VSS VSS VCC VCC _0394_ sky130_fd_sc_hd__nor2_1
X_3901_ net509 net98 net721 VSS VSS VCC VCC _1708_ sky130_fd_sc_hd__a21o_1
X_4881_ _2411_ _2414_ _2417_ net323 VSS VSS VCC VCC _2418_ sky130_fd_sc_hd__a31o_1
X_3832_ net510 _1655_ VSS VSS VCC VCC _1656_ sky130_fd_sc_hd__and2b_1
X_3763_ net654 net66 net395 VSS VSS VCC VCC _0032_ sky130_fd_sc_hd__mux2_1
X_2714_ _0686_ _0687_ net429 VSS VSS VCC VCC _0689_ sky130_fd_sc_hd__a21o_1
X_3694_ _0848_ _0907_ net608 VSS VSS VCC VCC _1573_ sky130_fd_sc_hd__a21boi_1
X_2645_ _0616_ _0617_ net429 VSS VSS VCC VCC _0620_ sky130_fd_sc_hd__a21o_1
Xoutput301 net301 VSS VSS VCC VCC o_wdata[2] sky130_fd_sc_hd__buf_2
Xoutput312 net312 VSS VSS VCC VCC o_wsel[1] sky130_fd_sc_hd__buf_2
X_5364_ clknet_leaf_68_i_clk _0391_ VSS VSS VCC VCC u_muldiv.mul\[43\] sky130_fd_sc_hd__dfxtp_1
X_2576_ net457 net537 _0460_ _0549_ VSS VSS VCC VCC _0551_ sky130_fd_sc_hd__o22ai_1
X_4315_ _1926_ _1931_ _1933_ _1942_ _1929_ VSS VSS VCC VCC _1943_ sky130_fd_sc_hd__a221o_1
X_5295_ clknet_4_9__leaf_i_clk _0323_ VSS VSS VCC VCC u_muldiv.dividend\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_4246_ _1873_ _1866_ _1871_ VSS VSS VCC VCC _1874_ sky130_fd_sc_hd__o21ai_2
X_4177_ u_muldiv.mul\[7\] u_muldiv.mul\[6\] net408 VSS VSS VCC VCC _0221_
+ sky130_fd_sc_hd__mux2_1
X_3128_ net654 net656 net658 net660 net637 net625 VSS VSS VCC VCC _1088_ sky130_fd_sc_hd__mux4_1
X_3059_ _1004_ _1022_ net735 VSS VSS VCC VCC _1023_ sky130_fd_sc_hd__a21oi_1
Xfanout550 u_muldiv.i_is_div VSS VSS VCC VCC net550 sky130_fd_sc_hd__buf_6
Xfanout561 net562 VSS VSS VCC VCC net561 sky130_fd_sc_hd__buf_4
Xfanout572 net215 VSS VSS VCC VCC net572 sky130_fd_sc_hd__clkbuf_4
Xfanout583 u_bits.i_op2\[26\] VSS VSS VCC VCC net583 sky130_fd_sc_hd__clkbuf_4
Xfanout594 u_bits.i_op2\[11\] VSS VSS VCC VCC net594 sky130_fd_sc_hd__clkbuf_16
X_4100_ u_bits.i_op2\[22\] u_bits.i_op2\[21\] _1779_ _1799_ VSS VSS VCC VCC
+ _1806_ sky130_fd_sc_hd__or4bb_4
X_5080_ clknet_leaf_125_i_clk _0113_ VSS VSS VCC VCC u_mux.i_group_mux sky130_fd_sc_hd__dfxtp_1
X_4031_ net597 _1750_ _1751_ VSS VSS VCC VCC _1752_ sky130_fd_sc_hd__o21ba_1
X_4933_ net461 _2434_ net474 VSS VSS VCC VCC _2435_ sky130_fd_sc_hd__mux2_1
X_4864_ u_muldiv.dividend\[29\] u_muldiv.dividend\[28\] u_muldiv.dividend\[27\] _2372_
+ VSS VSS VCC VCC _2402_ sky130_fd_sc_hd__or4_2
X_3815_ net596 net598 net549 VSS VSS VCC VCC _1643_ sky130_fd_sc_hd__mux2_1
X_4795_ net670 net672 _2316_ net370 net667 VSS VSS VCC VCC _2339_ sky130_fd_sc_hd__o311a_1
X_3746_ net693 net48 net395 VSS VSS VCC VCC _0015_ sky130_fd_sc_hd__mux2_1
X_3677_ u_muldiv.dividend\[18\] net420 net368 u_muldiv.o_div\[18\] net444 vssd1 vssd1
+ vccd1 vccd1 _1557_ sky130_fd_sc_hd__a221o_1
X_2628_ _0593_ _0602_ VSS VSS VCC VCC _0603_ sky130_fd_sc_hd__nor2_1
X_5347_ clknet_leaf_6_i_clk _0375_ VSS VSS VCC VCC u_muldiv.divisor\[30\]
+ sky130_fd_sc_hd__dfxtp_2
X_2559_ net542 u_muldiv.add_prev\[3\] VSS VSS VCC VCC _0534_ sky130_fd_sc_hd__and2_1
Xoutput186 net186 VSS VSS VCC VCC o_add[12] sky130_fd_sc_hd__buf_2
Xoutput197 net197 VSS VSS VCC VCC o_add[22] sky130_fd_sc_hd__buf_2
X_5278_ clknet_leaf_158_i_clk _0306_ VSS VSS VCC VCC u_muldiv.quotient_msk\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_4229_ u_muldiv.dividend\[1\] _0418_ VSS VSS VCC VCC _1857_ sky130_fd_sc_hd__or2_1
Xfanout380 net381 VSS VSS VCC VCC net380 sky130_fd_sc_hd__clkbuf_4
Xfanout391 net392 VSS VSS VCC VCC net391 sky130_fd_sc_hd__clkbuf_8
X_3600_ _1485_ _1484_ net356 _1198_ VSS VSS VCC VCC _1486_ sky130_fd_sc_hd__o22a_1
Xinput11 i_csr_data[14] VSS VSS VCC VCC net11 sky130_fd_sc_hd__buf_4
Xinput22 i_csr_data[24] VSS VSS VCC VCC net22 sky130_fd_sc_hd__buf_4
X_4580_ net460 net718 net715 net713 VSS VSS VCC VCC _2143_ sky130_fd_sc_hd__nor4_1
Xinput33 i_csr_data[5] VSS VSS VCC VCC net33 sky130_fd_sc_hd__buf_2
Xinput44 i_inst_jal_jalr VSS VSS VCC VCC net44 sky130_fd_sc_hd__buf_4
Xinput55 i_op1[19] VSS VSS VCC VCC net55 sky130_fd_sc_hd__clkbuf_1
X_3531_ net443 _1418_ _1421_ net734 VSS VSS VCC VCC _1422_ sky130_fd_sc_hd__a211o_1
Xinput66 i_op1[29] VSS VSS VCC VCC net66 sky130_fd_sc_hd__clkbuf_1
Xinput77 i_op2[0] VSS VSS VCC VCC net77 sky130_fd_sc_hd__buf_4
Xinput88 i_op2[1] VSS VSS VCC VCC net88 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput99 i_op2[2] VSS VSS VCC VCC net99 sky130_fd_sc_hd__buf_2
X_3462_ _1356_ net31 net733 VSS VSS VCC VCC _1357_ sky130_fd_sc_hd__mux2_2
X_5201_ clknet_leaf_154_i_clk _0233_ VSS VSS VCC VCC u_muldiv.mul\[18\] sky130_fd_sc_hd__dfxtp_1
X_3393_ _1289_ _1290_ _1288_ _1287_ VSS VSS VCC VCC _1291_ sky130_fd_sc_hd__o22ai_4
X_5132_ clknet_leaf_39_i_clk _0164_ VSS VSS VCC VCC u_muldiv.divisor\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_5063_ clknet_leaf_50_i_clk _0096_ VSS VSS VCC VCC net228 sky130_fd_sc_hd__dfxtp_4
X_4014_ net603 _1279_ net382 VSS VSS VCC VCC _1738_ sky130_fd_sc_hd__o21ai_1
X_4916_ u_muldiv.divisor\[23\] net476 net332 u_muldiv.divisor\[24\] vssd1 vssd1 vccd1
+ vccd1 _0368_ sky130_fd_sc_hd__a22o_1
X_4847_ _2378_ _2383_ _2386_ net315 VSS VSS VCC VCC _2387_ sky130_fd_sc_hd__o211a_1
X_4778_ net481 _2322_ _2323_ _2320_ VSS VSS VCC VCC _2324_ sky130_fd_sc_hd__a31o_1
X_3729_ _1596_ _1605_ net735 VSS VSS VCC VCC _1606_ sky130_fd_sc_hd__a21oi_4
X_2962_ u_muldiv.mul\[57\] net363 net357 u_muldiv.mul\[25\] VSS VSS VCC VCC
+ _0930_ sky130_fd_sc_hd__a22oi_1
X_4701_ _1905_ _2252_ VSS VSS VCC VCC _2253_ sky130_fd_sc_hd__xnor2_1
X_2893_ _0814_ _0851_ _0861_ _0864_ VSS VSS VCC VCC _0865_ sky130_fd_sc_hd__a31o_1
X_4632_ _1876_ _1879_ _1880_ _1844_ VSS VSS VCC VCC _2190_ sky130_fd_sc_hd__a22o_1
X_4563_ net498 _2126_ _2127_ _2121_ _2125_ VSS VSS VCC VCC _2128_ sky130_fd_sc_hd__a32o_1
X_3514_ u_muldiv.o_div\[6\] net366 net358 _1405_ VSS VSS VCC VCC _1406_ sky130_fd_sc_hd__a211o_1
X_4494_ u_muldiv.o_div\[28\] _2094_ VSS VSS VCC VCC _2095_ sky130_fd_sc_hd__or2_1
X_3445_ net696 net694 net692 net689 net646 net634 VSS VSS VCC VCC _1340_ sky130_fd_sc_hd__mux4_1
X_3376_ net460 net717 net715 net713 net643 net629 VSS VSS VCC VCC _1274_ sky130_fd_sc_hd__mux4_1
X_5115_ clknet_leaf_172_i_clk _0148_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[30\]
+ sky130_fd_sc_hd__dfxtp_2
X_5046_ clknet_leaf_51_i_clk _0079_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[4\]
+ sky130_fd_sc_hd__dfxtp_4
X_3230_ _1172_ _1176_ VSS VSS VCC VCC _1177_ sky130_fd_sc_hd__nand2_1
X_3161_ net612 _0777_ net347 VSS VSS VCC VCC _1119_ sky130_fd_sc_hd__o21ai_1
X_3092_ net560 _1053_ VSS VSS VCC VCC _1054_ sky130_fd_sc_hd__or2_1
X_3994_ u_muldiv.divisor\[31\] net477 net383 net640 VSS VSS VCC VCC _1723_
+ sky130_fd_sc_hd__a22o_1
X_2945_ _0900_ _0901_ _0912_ _0914_ _0895_ VSS VSS VCC VCC _0915_ sky130_fd_sc_hd__o2111ai_1
X_2876_ net712 net716 net717 net460 net644 net635 VSS VSS VCC VCC _0848_ sky130_fd_sc_hd__mux4_2
X_4615_ _0436_ _2172_ net373 _2174_ VSS VSS VCC VCC _2175_ sky130_fd_sc_hd__a31o_1
X_4546_ u_muldiv.divisor\[0\] _0440_ _2110_ _2111_ VSS VSS VCC VCC _2112_
+ sky130_fd_sc_hd__a31o_1
X_4477_ u_muldiv.o_div\[23\] _2074_ u_muldiv.o_div\[24\] VSS VSS VCC VCC _2082_
+ sky130_fd_sc_hd__o21ai_1
X_3428_ net610 _1323_ _0765_ _1321_ VSS VSS VCC VCC _1324_ sky130_fd_sc_hd__o211a_1
X_3359_ u_wr_mux.i_reg_data2\[13\] _0764_ _1263_ VSS VSS VCC VCC net300 sky130_fd_sc_hd__a21o_1
X_5029_ clknet_leaf_52_i_clk _0062_ VSS VSS VCC VCC u_bits.i_op2\[18\] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_1_i_clk clknet_4_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2730_ _0700_ _0703_ _0702_ VSS VSS VCC VCC _0705_ sky130_fd_sc_hd__o21ai_1
X_2661_ _0584_ _0603_ _0634_ VSS VSS VCC VCC _0636_ sky130_fd_sc_hd__nand3_4
X_4400_ _0452_ _2019_ VSS VSS VCC VCC _2021_ sky130_fd_sc_hd__or2_1
X_5380_ clknet_4_3__leaf_i_clk _0407_ VSS VSS VCC VCC u_muldiv.mul\[59\] sky130_fd_sc_hd__dfxtp_1
X_2592_ net718 u_muldiv.add_prev\[1\] net537 VSS VSS VCC VCC _0567_ sky130_fd_sc_hd__mux2_1
X_4331_ _1950_ _1953_ _1957_ _1958_ _1951_ VSS VSS VCC VCC _1959_ sky130_fd_sc_hd__o311a_1
X_4262_ _0416_ u_muldiv.dividend\[11\] _1885_ VSS VSS VCC VCC _1890_ sky130_fd_sc_hd__o21ai_1
X_3213_ _0568_ _0578_ _0562_ VSS VSS VCC VCC _1164_ sky130_fd_sc_hd__a21o_1
X_4193_ u_muldiv.mul\[23\] u_muldiv.mul\[22\] net405 VSS VSS VCC VCC _0237_
+ sky130_fd_sc_hd__mux2_1
X_3144_ net427 _1102_ VSS VSS VCC VCC _1103_ sky130_fd_sc_hd__xor2_1
X_3075_ u_muldiv.dividend\[28\] net419 net364 u_muldiv.o_div\[28\] net442 vssd1 vssd1
+ vccd1 vccd1 _1037_ sky130_fd_sc_hd__a221o_1
X_3977_ u_wr_mux.i_reg_data2\[21\] net157 net395 VSS VSS VCC VCC _0139_ sky130_fd_sc_hd__mux2_1
X_2928_ net711 net712 net715 net718 net649 net634 VSS VSS VCC VCC _0898_ sky130_fd_sc_hd__mux4_1
X_2859_ _0830_ _0831_ VSS VSS VCC VCC _0832_ sky130_fd_sc_hd__xnor2_4
X_4529_ u_muldiv.quotient_msk\[17\] net491 net340 u_muldiv.quotient_msk\[18\] vssd1
+ vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__a22o_1
Xfanout710 net711 VSS VSS VCC VCC net710 sky130_fd_sc_hd__buf_6
Xfanout721 net722 VSS VSS VCC VCC net721 sky130_fd_sc_hd__buf_4
Xfanout732 _0424_ VSS VSS VCC VCC net732 sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_164_i_clk clknet_4_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_164_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_102_i_clk clknet_4_12__leaf_i_clk VSS VSS VCC VCC clknet_leaf_102_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput9 i_csr_data[12] VSS VSS VCC VCC net9 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_117_i_clk clknet_4_11__leaf_i_clk VSS VSS VCC VCC clknet_leaf_117_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3900_ net509 _1706_ VSS VSS VCC VCC _1707_ sky130_fd_sc_hd__and2b_1
X_4880_ net652 _2415_ _2416_ VSS VSS VCC VCC _2417_ sky130_fd_sc_hd__a21o_1
X_3831_ net592 net594 net550 VSS VSS VCC VCC _1655_ sky130_fd_sc_hd__mux2_1
X_3762_ net657 net65 net390 VSS VSS VCC VCC _0031_ sky130_fd_sc_hd__mux2_1
X_2713_ _0686_ _0687_ net429 VSS VSS VCC VCC _0688_ sky130_fd_sc_hd__a21oi_1
X_3693_ net608 _1338_ net328 VSS VSS VCC VCC _1572_ sky130_fd_sc_hd__o21ai_1
X_2644_ _0616_ _0617_ net431 VSS VSS VCC VCC _0619_ sky130_fd_sc_hd__a21o_1
Xoutput302 net302 VSS VSS VCC VCC o_wdata[30] sky130_fd_sc_hd__buf_2
Xoutput313 net313 VSS VSS VCC VCC o_wsel[2] sky130_fd_sc_hd__buf_2
X_5363_ clknet_leaf_77_i_clk _0390_ VSS VSS VCC VCC u_muldiv.mul\[42\] sky130_fd_sc_hd__dfxtp_2
X_2575_ net646 net551 net716 net537 net423 VSS VSS VCC VCC _0550_ sky130_fd_sc_hd__o2111ai_1
X_4314_ _1938_ _1934_ _1939_ VSS VSS VCC VCC _1942_ sky130_fd_sc_hd__a21o_1
X_5294_ clknet_4_11__leaf_i_clk _0322_ VSS VSS VCC VCC u_muldiv.dividend\[9\]
+ sky130_fd_sc_hd__dfxtp_4
X_4245_ _1867_ _1872_ VSS VSS VCC VCC _1873_ sky130_fd_sc_hd__nand2_1
X_4176_ u_muldiv.mul\[6\] u_muldiv.mul\[5\] net403 VSS VSS VCC VCC _0220_
+ sky130_fd_sc_hd__mux2_1
X_3127_ net453 _0944_ _1086_ VSS VSS VCC VCC _1087_ sky130_fd_sc_hd__o21ai_1
X_3058_ net355 _1000_ _1001_ _1021_ net532 VSS VSS VCC VCC _1022_ sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_81_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_81_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_96_i_clk clknet_4_14__leaf_i_clk VSS VSS VCC VCC clknet_leaf_96_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout540 net543 VSS VSS VCC VCC net540 sky130_fd_sc_hd__buf_6
Xfanout551 net553 VSS VSS VCC VCC net551 sky130_fd_sc_hd__buf_4
Xfanout562 net563 VSS VSS VCC VCC net562 sky130_fd_sc_hd__buf_6
Xfanout573 net215 VSS VSS VCC VCC net573 sky130_fd_sc_hd__buf_4
Xfanout584 u_bits.i_op2\[25\] VSS VSS VCC VCC net584 sky130_fd_sc_hd__buf_4
Xfanout595 u_bits.i_op2\[10\] VSS VSS VCC VCC net595 sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_34_i_clk clknet_4_4__leaf_i_clk VSS VSS VCC VCC clknet_leaf_34_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_49_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_49_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4030_ _1749_ net379 net597 net329 VSS VSS VCC VCC _1751_ sky130_fd_sc_hd__a31o_1
X_4932_ _1859_ _2433_ VSS VSS VCC VCC _2434_ sky130_fd_sc_hd__nand2_1
X_4863_ u_muldiv.dividend\[28\] u_muldiv.dividend\[27\] _2372_ u_muldiv.dividend\[29\]
+ VSS VSS VCC VCC _2401_ sky130_fd_sc_hd__o31a_1
X_3814_ net598 net725 _1642_ _1641_ VSS VSS VCC VCC _0051_ sky130_fd_sc_hd__o22a_1
X_4794_ net670 net672 _2316_ VSS VSS VCC VCC _2338_ sky130_fd_sc_hd__or3_4
X_3745_ net695 net47 net393 VSS VSS VCC VCC _0014_ sky130_fd_sc_hd__mux2_1
X_3676_ net731 _1555_ _1556_ net578 VSS VSS VCC VCC net253 sky130_fd_sc_hd__a211oi_4
X_2627_ _0600_ _0601_ VSS VSS VCC VCC _0602_ sky130_fd_sc_hd__nand2_1
X_2558_ _0525_ _0530_ _0529_ _0510_ VSS VSS VCC VCC _0533_ sky130_fd_sc_hd__nor4_2
X_5346_ clknet_leaf_6_i_clk _0374_ VSS VSS VCC VCC u_muldiv.divisor\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput187 net187 VSS VSS VCC VCC o_add[13] sky130_fd_sc_hd__buf_2
Xoutput198 net198 VSS VSS VCC VCC o_add[23] sky130_fd_sc_hd__buf_2
X_2489_ net641 net549 net534 net424 VSS VSS VCC VCC _0464_ sky130_fd_sc_hd__o211a_2
X_5277_ clknet_leaf_161_i_clk _0305_ VSS VSS VCC VCC u_muldiv.quotient_msk\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_4228_ _0417_ net463 VSS VSS VCC VCC _1856_ sky130_fd_sc_hd__nand2_1
X_4159_ net552 net500 net195 VSS VSS VCC VCC _0203_ sky130_fd_sc_hd__o21a_1
Xfanout370 net371 VSS VSS VCC VCC net370 sky130_fd_sc_hd__buf_2
Xfanout381 net382 VSS VSS VCC VCC net381 sky130_fd_sc_hd__clkbuf_4
Xfanout392 _1610_ VSS VSS VCC VCC net392 sky130_fd_sc_hd__clkbuf_4
Xinput12 i_csr_data[15] VSS VSS VCC VCC net12 sky130_fd_sc_hd__buf_4
Xinput23 i_csr_data[25] VSS VSS VCC VCC net23 sky130_fd_sc_hd__clkbuf_4
Xinput34 i_csr_data[6] VSS VSS VCC VCC net34 sky130_fd_sc_hd__clkbuf_4
Xinput45 i_op1[0] VSS VSS VCC VCC net45 sky130_fd_sc_hd__clkbuf_2
X_3530_ net559 u_muldiv.mul\[7\] net413 net528 _1420_ VSS VSS VCC VCC _1421_
+ sky130_fd_sc_hd__o311a_1
Xinput56 i_op1[1] VSS VSS VCC VCC net56 sky130_fd_sc_hd__clkbuf_1
Xinput67 i_op1[2] VSS VSS VCC VCC net67 sky130_fd_sc_hd__clkbuf_1
Xinput78 i_op2[10] VSS VSS VCC VCC net78 sky130_fd_sc_hd__clkbuf_1
Xinput89 i_op2[20] VSS VSS VCC VCC net89 sky130_fd_sc_hd__clkbuf_1
X_3461_ _1355_ _1354_ _1352_ net447 VSS VSS VCC VCC _1356_ sky130_fd_sc_hd__a22o_2
X_5200_ clknet_leaf_154_i_clk _0232_ VSS VSS VCC VCC u_muldiv.mul\[17\] sky130_fd_sc_hd__dfxtp_1
X_3392_ u_muldiv.dividend\[0\] net420 net367 u_muldiv.o_div\[0\] net447 vssd1 vssd1
+ vccd1 vccd1 _1290_ sky130_fd_sc_hd__a221o_2
X_5131_ clknet_4_6__leaf_i_clk _0163_ VSS VSS VCC VCC u_muldiv.divisor\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_5062_ clknet_leaf_133_i_clk _0095_ VSS VSS VCC VCC net227 sky130_fd_sc_hd__dfxtp_1
X_4013_ net603 u_bits.i_op2\[0\] net636 _0908_ VSS VSS VCC VCC _1737_ sky130_fd_sc_hd__or4_1
X_4915_ u_muldiv.divisor\[22\] net480 net334 u_muldiv.divisor\[23\] vssd1 vssd1 vccd1
+ vccd1 _0367_ sky130_fd_sc_hd__a22o_1
X_4846_ u_muldiv.dividend\[27\] _2372_ _2385_ VSS VSS VCC VCC _2386_ sky130_fd_sc_hd__o21ai_1
X_4777_ u_muldiv.dividend\[20\] u_muldiv.dividend\[19\] _2284_ u_muldiv.dividend\[21\]
+ VSS VSS VCC VCC _2323_ sky130_fd_sc_hd__o31ai_1
X_3728_ net520 _1604_ net356 _1210_ net442 VSS VSS VCC VCC _1605_ sky130_fd_sc_hd__o221ai_4
X_3659_ _1539_ _1540_ VSS VSS VCC VCC _1541_ sky130_fd_sc_hd__nor2_1
X_5329_ clknet_leaf_137_i_clk _0357_ VSS VSS VCC VCC u_muldiv.divisor\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_2961_ u_muldiv.dividend\[25\] net419 net364 u_muldiv.o_div\[25\] vssd1 vssd1 vccd1
+ vccd1 _0929_ sky130_fd_sc_hd__a22oi_2
X_4700_ _0414_ u_muldiv.dividend\[14\] _2245_ VSS VSS VCC VCC _2252_ sky130_fd_sc_hd__a21oi_1
X_2892_ net669 net586 net411 _0844_ _0863_ VSS VSS VCC VCC _0864_ sky130_fd_sc_hd__a311o_1
X_4631_ u_muldiv.dividend\[8\] net324 net375 _2189_ VSS VSS VCC VCC _0321_
+ sky130_fd_sc_hd__a31o_1
X_4562_ u_muldiv.dividend\[0\] net464 net463 VSS VSS VCC VCC _2127_ sky130_fd_sc_hd__o21ai_1
X_3513_ net567 net556 u_muldiv.dividend\[6\] u_muldiv.mul\[38\] net361 vssd1 vssd1
+ vccd1 vccd1 _1405_ sky130_fd_sc_hd__a32o_1
X_4493_ u_muldiv.o_div\[25\] u_muldiv.o_div\[26\] u_muldiv.o_div\[27\] _2081_ vssd1
+ vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__or4_2
X_3444_ net687 net685 u_bits.i_op1\[17\] net681 net646 net634 VSS VSS VCC VCC
+ _1339_ sky130_fd_sc_hd__mux4_1
X_3375_ net710 net708 net706 net704 net643 net628 VSS VSS VCC VCC _1273_ sky130_fd_sc_hd__mux4_1
X_5114_ clknet_leaf_35_i_clk _0147_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_5045_ clknet_leaf_91_i_clk _0078_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[3\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_4_7__f_i_clk clknet_2_1_0_i_clk VSS VSS VCC VCC clknet_4_7__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4829_ _2368_ net369 net660 net465 VSS VSS VCC VCC _2370_ sky130_fd_sc_hd__a31oi_1
X_3160_ net612 _0777_ _0890_ VSS VSS VCC VCC _1118_ sky130_fd_sc_hd__o21a_1
Xhold1 u_muldiv.mul\[8\] VSS VSS VCC VCC net736 sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ net657 u_bits.i_op2\[28\] VSS VSS VCC VCC _1053_ sky130_fd_sc_hd__nand2_1
X_3993_ _0413_ net436 VSS VSS VCC VCC _1722_ sky130_fd_sc_hd__nand2_1
X_2944_ net664 net585 _0913_ net348 VSS VSS VCC VCC _0914_ sky130_fd_sc_hd__o211ai_1
X_2875_ net458 net717 _0846_ VSS VSS VCC VCC _0847_ sky130_fd_sc_hd__a21boi_2
X_4614_ _2173_ net704 net472 VSS VSS VCC VCC _2174_ sky130_fd_sc_hd__a21o_1
X_4545_ _1857_ _1858_ _1859_ net459 VSS VSS VCC VCC _2111_ sky130_fd_sc_hd__a31o_1
X_4476_ u_muldiv.o_div\[23\] u_muldiv.o_div\[24\] _2074_ VSS VSS VCC VCC _2081_
+ sky130_fd_sc_hd__or3_4
X_3427_ _1316_ _1317_ _1322_ _1318_ net621 net451 VSS VSS VCC VCC _1323_ sky130_fd_sc_hd__mux4_1
X_3358_ net562 u_wr_mux.i_reg_data2\[29\] net416 net306 VSS VSS VCC VCC _1263_
+ sky130_fd_sc_hd__a22o_1
X_3289_ _0530_ _0743_ _0525_ VSS VSS VCC VCC _1220_ sky130_fd_sc_hd__o21ba_1
X_5028_ clknet_4_5__leaf_i_clk _0061_ VSS VSS VCC VCC u_bits.i_op2\[17\] sky130_fd_sc_hd__dfxtp_4
X_2660_ _0632_ _0633_ _0627_ VSS VSS VCC VCC _0635_ sky130_fd_sc_hd__o21ai_2
X_2591_ _0563_ _0564_ net431 VSS VSS VCC VCC _0566_ sky130_fd_sc_hd__a21o_1
X_4330_ u_muldiv.divisor\[27\] _0448_ _1948_ VSS VSS VCC VCC _1958_ sky130_fd_sc_hd__a21o_1
X_4261_ _1885_ _1886_ _1888_ VSS VSS VCC VCC _1889_ sky130_fd_sc_hd__or3_1
X_3212_ _1162_ _1163_ VSS VSS VCC VCC net208 sky130_fd_sc_hd__nand2_4
X_4192_ u_muldiv.mul\[22\] u_muldiv.mul\[21\] net405 VSS VSS VCC VCC _0236_
+ sky130_fd_sc_hd__mux2_1
X_3143_ net445 net580 _0464_ net653 VSS VSS VCC VCC _1102_ sky130_fd_sc_hd__a22o_1
X_3074_ _1030_ _1036_ VSS VSS VCC VCC net203 sky130_fd_sc_hd__xnor2_4
X_3976_ u_wr_mux.i_reg_data2\[20\] net156 net392 VSS VSS VCC VCC _0138_ sky130_fd_sc_hd__mux2_1
X_2927_ net454 net613 VSS VSS VCC VCC _0897_ sky130_fd_sc_hd__nand2_1
X_2858_ _0468_ _0471_ _0750_ _0473_ VSS VSS VCC VCC _0831_ sky130_fd_sc_hd__a22oi_4
X_2789_ net417 net441 net522 VSS VSS VCC VCC _0763_ sky130_fd_sc_hd__a21o_1
X_4528_ u_muldiv.quotient_msk\[16\] net491 net338 u_muldiv.quotient_msk\[17\] vssd1
+ vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__a22o_1
Xfanout700 u_bits.i_op1\[9\] VSS VSS VCC VCC net700 sky130_fd_sc_hd__clkbuf_16
X_4459_ u_muldiv.quotient_msk\[20\] u_muldiv.o_div\[20\] net469 net437 vssd1 vssd1
+ vccd1 vccd1 _2068_ sky130_fd_sc_hd__o211a_1
Xfanout711 u_bits.i_op1\[4\] VSS VSS VCC VCC net711 sky130_fd_sc_hd__buf_6
Xfanout722 _1609_ VSS VSS VCC VCC net722 sky130_fd_sc_hd__clkbuf_4
Xfanout733 net38 VSS VSS VCC VCC net733 sky130_fd_sc_hd__buf_6
X_3830_ net594 net725 _1654_ _1653_ VSS VSS VCC VCC _0055_ sky130_fd_sc_hd__o22a_1
X_3761_ net659 net64 net389 VSS VSS VCC VCC _0030_ sky130_fd_sc_hd__mux2_1
X_2712_ net449 net595 VSS VSS VCC VCC _0687_ sky130_fd_sc_hd__nand2_1
X_3692_ u_muldiv.mul\[51\] net361 net360 u_muldiv.mul\[19\] _1570_ vssd1 vssd1 vccd1
+ vccd1 _1571_ sky130_fd_sc_hd__a221oi_1
X_2643_ _0616_ _0617_ net431 VSS VSS VCC VCC _0618_ sky130_fd_sc_hd__nand3_1
Xoutput303 net303 VSS VSS VCC VCC o_wdata[31] sky130_fd_sc_hd__buf_2
Xoutput314 net314 VSS VSS VCC VCC o_wsel[3] sky130_fd_sc_hd__buf_2
X_5362_ clknet_leaf_76_i_clk _0389_ VSS VSS VCC VCC u_muldiv.mul\[41\] sky130_fd_sc_hd__dfxtp_2
X_2574_ net646 net551 net716 net538 VSS VSS VCC VCC _0549_ sky130_fd_sc_hd__o211ai_4
X_4313_ _1926_ _1940_ _1927_ _1932_ VSS VSS VCC VCC _1941_ sky130_fd_sc_hd__or4b_1
X_5293_ clknet_4_11__leaf_i_clk _0321_ VSS VSS VCC VCC u_muldiv.dividend\[8\]
+ sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_0_i_clk clknet_4_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4244_ _1845_ _1846_ VSS VSS VCC VCC _1872_ sky130_fd_sc_hd__and2_1
X_4175_ u_muldiv.mul\[5\] u_muldiv.mul\[4\] net403 VSS VSS VCC VCC _0219_
+ sky130_fd_sc_hd__mux2_1
X_3126_ net619 _0947_ VSS VSS VCC VCC _1086_ sky130_fd_sc_hd__or2_1
X_3057_ _1007_ _1020_ _0422_ VSS VSS VCC VCC _1021_ sky130_fd_sc_hd__o21a_1
X_3959_ net304 net169 net387 VSS VSS VCC VCC _0121_ sky130_fd_sc_hd__mux2_1
Xfanout530 net544 VSS VSS VCC VCC net530 sky130_fd_sc_hd__buf_4
Xfanout541 net543 VSS VSS VCC VCC net541 sky130_fd_sc_hd__clkbuf_4
Xfanout552 net553 VSS VSS VCC VCC net552 sky130_fd_sc_hd__buf_6
Xfanout563 net216 VSS VSS VCC VCC net563 sky130_fd_sc_hd__clkbuf_16
Xfanout574 net575 VSS VSS VCC VCC net574 sky130_fd_sc_hd__buf_6
Xfanout585 u_bits.i_op2\[24\] VSS VSS VCC VCC net585 sky130_fd_sc_hd__buf_4
Xfanout596 u_bits.i_op2\[9\] VSS VSS VCC VCC net596 sky130_fd_sc_hd__buf_6
X_4931_ u_muldiv.divisor\[0\] _0440_ VSS VSS VCC VCC _2433_ sky130_fd_sc_hd__or2_1
X_4862_ _1962_ _1963_ _2398_ _1720_ VSS VSS VCC VCC _2400_ sky130_fd_sc_hd__a31o_1
X_3813_ net505 net106 net719 VSS VSS VCC VCC _1642_ sky130_fd_sc_hd__a21o_1
X_4793_ _1930_ _1931_ _2335_ _2336_ VSS VSS VCC VCC _2337_ sky130_fd_sc_hd__a31o_1
X_3744_ net698 net46 net399 VSS VSS VCC VCC _0013_ sky130_fd_sc_hd__mux2_1
X_3675_ net14 net732 VSS VSS VCC VCC _1556_ sky130_fd_sc_hd__nor2_2
X_2626_ _0596_ _0597_ _0598_ VSS VSS VCC VCC _0601_ sky130_fd_sc_hd__nand3_4
X_5345_ clknet_leaf_3_i_clk _0373_ VSS VSS VCC VCC u_muldiv.divisor\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_2557_ _0531_ _0519_ _0518_ VSS VSS VCC VCC _0532_ sky130_fd_sc_hd__and3_1
Xoutput188 net188 VSS VSS VCC VCC o_add[14] sky130_fd_sc_hd__buf_2
X_5276_ clknet_leaf_153_i_clk _0304_ VSS VSS VCC VCC u_muldiv.quotient_msk\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput199 net199 VSS VSS VCC VCC o_add[24] sky130_fd_sc_hd__buf_2
X_2488_ net551 _0419_ _0462_ VSS VSS VCC VCC _0463_ sky130_fd_sc_hd__o21ai_4
X_4227_ _0442_ u_muldiv.divisor\[2\] VSS VSS VCC VCC _1855_ sky130_fd_sc_hd__nand2_1
X_4158_ net553 u_muldiv.i_on_wait net193 VSS VSS VCC VCC _0202_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_163_i_clk clknet_4_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_163_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3109_ _1030_ _1035_ _1029_ VSS VSS VCC VCC _1070_ sky130_fd_sc_hd__o21ai_1
X_4089_ u_bits.i_op2\[20\] _1796_ _1797_ VSS VSS VCC VCC _1798_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_178_i_clk clknet_4_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_178_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_116_i_clk clknet_4_11__leaf_i_clk VSS VSS VCC VCC clknet_leaf_116_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout360 _0760_ VSS VSS VCC VCC net360 sky130_fd_sc_hd__buf_6
Xfanout371 _2113_ VSS VSS VCC VCC net371 sky130_fd_sc_hd__clkbuf_4
Xfanout382 _1724_ VSS VSS VCC VCC net382 sky130_fd_sc_hd__clkbuf_4
Xfanout393 net394 VSS VSS VCC VCC net393 sky130_fd_sc_hd__buf_4
Xinput13 i_csr_data[16] VSS VSS VCC VCC net13 sky130_fd_sc_hd__buf_6
Xinput24 i_csr_data[26] VSS VSS VCC VCC net24 sky130_fd_sc_hd__clkbuf_2
Xinput35 i_csr_data[7] VSS VSS VCC VCC net35 sky130_fd_sc_hd__buf_6
Xinput46 i_op1[10] VSS VSS VCC VCC net46 sky130_fd_sc_hd__clkbuf_1
Xinput57 i_op1[20] VSS VSS VCC VCC net57 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput68 i_op1[30] VSS VSS VCC VCC net68 sky130_fd_sc_hd__clkbuf_1
Xinput79 i_op2[11] VSS VSS VCC VCC net79 sky130_fd_sc_hd__clkbuf_4
X_3460_ net557 u_muldiv.mul\[3\] net414 net529 VSS VSS VCC VCC _1355_ sky130_fd_sc_hd__o31a_1
X_3391_ u_muldiv.mul\[32\] net361 net359 u_muldiv.mul\[0\] VSS VSS VCC VCC
+ _1289_ sky130_fd_sc_hd__a22o_1
X_5130_ clknet_leaf_37_i_clk _0162_ VSS VSS VCC VCC u_muldiv.divisor\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_5061_ clknet_leaf_166_i_clk _0094_ VSS VSS VCC VCC net226 sky130_fd_sc_hd__dfxtp_2
X_4012_ u_muldiv.divisor\[35\] net478 net333 u_muldiv.divisor\[36\] _1736_ vssd1 vssd1
+ vccd1 vccd1 _0155_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_95_i_clk clknet_4_14__leaf_i_clk VSS VSS VCC VCC clknet_leaf_95_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4914_ u_muldiv.divisor\[21\] net480 net334 u_muldiv.divisor\[22\] vssd1 vssd1 vccd1
+ vccd1 _0366_ sky130_fd_sc_hd__a22o_1
X_4845_ _2372_ u_muldiv.dividend\[27\] net433 VSS VSS VCC VCC _2385_ sky130_fd_sc_hd__a21oi_1
X_4776_ _2280_ _2321_ _0450_ VSS VSS VCC VCC _2322_ sky130_fd_sc_hd__nand3_2
X_3727_ _0814_ _1603_ _1600_ _1597_ VSS VSS VCC VCC _1604_ sky130_fd_sc_hd__a211oi_2
X_3658_ u_bits.i_op2\[16\] u_bits.i_op1\[16\] net412 _1535_ _1537_ vssd1 vssd1 vccd1
+ vccd1 _1540_ sky130_fd_sc_hd__a311o_1
X_2609_ _0582_ _0583_ VSS VSS VCC VCC _0584_ sky130_fd_sc_hd__nand2_2
X_3589_ net556 u_muldiv.mul\[11\] net413 net528 VSS VSS VCC VCC _1476_ sky130_fd_sc_hd__o31a_1
X_5328_ clknet_4_8__leaf_i_clk _0356_ VSS VSS VCC VCC u_muldiv.divisor\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_48_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_48_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5259_ clknet_leaf_116_i_clk _0287_ VSS VSS VCC VCC u_muldiv.quotient_msk\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2960_ _0928_ VSS VSS VCC VCC net200 sky130_fd_sc_hd__clkinv_2
X_2891_ net669 u_bits.i_op2\[23\] _0862_ net348 VSS VSS VCC VCC _0863_ sky130_fd_sc_hd__o211a_1
X_4630_ _2188_ _2187_ _2182_ net318 VSS VSS VCC VCC _2189_ sky130_fd_sc_hd__o211a_1
X_4561_ u_muldiv.dividend\[0\] net464 net463 VSS VSS VCC VCC _2126_ sky130_fd_sc_hd__or3_1
X_3512_ _1403_ _1402_ net211 net354 VSS VSS VCC VCC _1404_ sky130_fd_sc_hd__a2bb2o_1
X_4492_ net323 _2091_ _2093_ VSS VSS VCC VCC _0278_ sky130_fd_sc_hd__o21a_1
X_3443_ _0836_ _0841_ _1337_ _0837_ net623 net452 VSS VSS VCC VCC _1338_ sky130_fd_sc_hd__mux4_2
X_3374_ _0891_ _0892_ _1270_ _1271_ net619 net450 VSS VSS VCC VCC _1272_ sky130_fd_sc_hd__mux4_2
X_5113_ clknet_leaf_94_i_clk _0146_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[28\]
+ sky130_fd_sc_hd__dfxtp_2
X_5044_ clknet_leaf_129_i_clk _0077_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4828_ net662 net369 _2358_ net660 VSS VSS VCC VCC _2369_ sky130_fd_sc_hd__a211o_1
X_4759_ _2304_ _2305_ net481 VSS VSS VCC VCC _2306_ sky130_fd_sc_hd__o21ai_1
Xhold2 u_muldiv.divisor\[43\] VSS VSS VCC VCC net737 sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ net611 _1049_ _1051_ VSS VSS VCC VCC _1052_ sky130_fd_sc_hd__a21oi_1
X_3992_ net465 net475 VSS VSS VCC VCC _1721_ sky130_fd_sc_hd__nor2_1
X_2943_ net560 net585 net665 VSS VSS VCC VCC _0913_ sky130_fd_sc_hd__nand3b_1
X_2874_ net644 net460 VSS VSS VCC VCC _0846_ sky130_fd_sc_hd__nand2_1
X_4613_ _2143_ _2171_ _0435_ _2114_ VSS VSS VCC VCC _2173_ sky130_fd_sc_hd__a31o_1
X_4544_ _1857_ _1858_ VSS VSS VCC VCC _2110_ sky130_fd_sc_hd__nand2_1
X_4475_ net317 _2078_ _2080_ VSS VSS VCC VCC _0274_ sky130_fd_sc_hd__a21oi_1
X_3426_ net715 net712 net710 net708 net645 net632 VSS VSS VCC VCC _1322_ sky130_fd_sc_hd__mux4_1
X_3357_ u_wr_mux.i_reg_data2\[12\] _0764_ _1262_ VSS VSS VCC VCC net299 sky130_fd_sc_hd__a21o_2
X_3288_ _1219_ VSS VSS VCC VCC net190 sky130_fd_sc_hd__inv_2
X_5027_ clknet_leaf_23_i_clk _0060_ VSS VSS VCC VCC u_bits.i_op2\[16\] sky130_fd_sc_hd__dfxtp_2
X_2590_ _0563_ _0564_ net431 VSS VSS VCC VCC _0565_ sky130_fd_sc_hd__nand3_1
X_4260_ u_muldiv.divisor\[11\] u_muldiv.dividend\[11\] VSS VSS VCC VCC _1888_
+ sky130_fd_sc_hd__xor2_1
X_3211_ _0560_ _0579_ _0581_ VSS VSS VCC VCC _1163_ sky130_fd_sc_hd__a21o_1
X_4191_ u_muldiv.mul\[21\] u_muldiv.mul\[20\] net404 VSS VSS VCC VCC _0235_
+ sky130_fd_sc_hd__mux2_1
X_3142_ _1036_ _1098_ _1100_ VSS VSS VCC VCC _1101_ sky130_fd_sc_hd__a21boi_2
X_3073_ _1032_ _0887_ _1034_ VSS VSS VCC VCC _1036_ sky130_fd_sc_hd__o21bai_4
X_3975_ u_wr_mux.i_reg_data2\[19\] net154 net399 VSS VSS VCC VCC _0137_ sky130_fd_sc_hd__mux2_1
X_2926_ net628 _0791_ VSS VSS VCC VCC _0896_ sky130_fd_sc_hd__nor2_1
X_2857_ _0828_ _0829_ VSS VSS VCC VCC _0830_ sky130_fd_sc_hd__nand2_2
X_2788_ net566 net556 net572 _0422_ VSS VSS VCC VCC _0762_ sky130_fd_sc_hd__o31a_2
X_4527_ u_muldiv.quotient_msk\[15\] net490 net338 u_muldiv.quotient_msk\[16\] vssd1
+ vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__a22o_1
X_4458_ u_muldiv.o_div\[18\] u_muldiv.o_div\[19\] _2058_ u_muldiv.o_div\[20\] vssd1
+ vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__o31ai_1
Xfanout701 net702 VSS VSS VCC VCC net701 sky130_fd_sc_hd__buf_4
Xfanout712 net713 VSS VSS VCC VCC net712 sky130_fd_sc_hd__buf_4
Xfanout723 net724 VSS VSS VCC VCC net723 sky130_fd_sc_hd__clkbuf_4
X_3409_ net632 net717 _1305_ net350 VSS VSS VCC VCC _1306_ sky130_fd_sc_hd__o211a_1
X_4389_ u_muldiv.o_div\[4\] u_muldiv.o_div\[5\] u_muldiv.o_div\[6\] _2005_ vssd1 vssd1
+ vccd1 vccd1 _2012_ sky130_fd_sc_hd__nor4_2
Xfanout734 net735 VSS VSS VCC VCC net734 sky130_fd_sc_hd__buf_2
X_3760_ u_bits.i_op1\[26\] net63 net393 VSS VSS VCC VCC _0029_ sky130_fd_sc_hd__mux2_1
X_2711_ net648 net554 net698 net540 net426 VSS VSS VCC VCC _0686_ sky130_fd_sc_hd__o2111ai_4
X_3691_ u_muldiv.dividend\[19\] net420 net368 u_muldiv.o_div\[19\] vssd1 vssd1 vccd1
+ vccd1 _1570_ sky130_fd_sc_hd__a22o_1
X_2642_ net447 u_bits.i_op2\[6\] VSS VSS VCC VCC _0617_ sky130_fd_sc_hd__nand2_1
X_5361_ clknet_leaf_75_i_clk _0388_ VSS VSS VCC VCC u_muldiv.mul\[40\] sky130_fd_sc_hd__dfxtp_2
Xoutput304 net304 VSS VSS VCC VCC o_wdata[3] sky130_fd_sc_hd__buf_2
X_2573_ net447 u_bits.i_op2\[2\] VSS VSS VCC VCC _0548_ sky130_fd_sc_hd__nand2_1
X_4312_ _1934_ _1935_ _1937_ _1939_ VSS VSS VCC VCC _1940_ sky130_fd_sc_hd__or4_1
X_5292_ clknet_leaf_122_i_clk _0320_ VSS VSS VCC VCC u_muldiv.dividend\[7\]
+ sky130_fd_sc_hd__dfxtp_4
X_4243_ _1846_ _1870_ VSS VSS VCC VCC _1871_ sky130_fd_sc_hd__and2_1
X_4174_ u_muldiv.mul\[4\] u_muldiv.mul\[3\] net403 VSS VSS VCC VCC _0218_
+ sky130_fd_sc_hd__mux2_1
X_3125_ net655 net581 net348 _1084_ VSS VSS VCC VCC _1085_ sky130_fd_sc_hd__o211a_1
X_3056_ _1011_ _0814_ net603 _1019_ _1016_ VSS VSS VCC VCC _1020_ sky130_fd_sc_hd__a311o_1
X_3958_ net301 net166 net391 VSS VSS VCC VCC _0120_ sky130_fd_sc_hd__mux2_1
X_2909_ _0533_ _0879_ VSS VSS VCC VCC _0880_ sky130_fd_sc_hd__nand2_2
X_3889_ net501 net95 net720 VSS VSS VCC VCC _1699_ sky130_fd_sc_hd__a21o_1
Xfanout520 net521 VSS VSS VCC VCC net520 sky130_fd_sc_hd__clkbuf_8
Xfanout531 net532 VSS VSS VCC VCC net531 sky130_fd_sc_hd__buf_4
Xfanout542 net543 VSS VSS VCC VCC net542 sky130_fd_sc_hd__buf_6
Xfanout553 net554 VSS VSS VCC VCC net553 sky130_fd_sc_hd__buf_4
Xfanout564 net569 VSS VSS VCC VCC net564 sky130_fd_sc_hd__buf_4
Xfanout575 net576 VSS VSS VCC VCC net575 sky130_fd_sc_hd__buf_6
Xfanout586 u_bits.i_op2\[23\] VSS VSS VCC VCC net586 sky130_fd_sc_hd__buf_4
Xfanout597 u_bits.i_op2\[8\] VSS VSS VCC VCC net597 sky130_fd_sc_hd__buf_6
X_4930_ net473 net497 _2432_ VSS VSS VCC VCC _0377_ sky130_fd_sc_hd__o21a_1
X_4861_ _1962_ _1963_ _2398_ VSS VSS VCC VCC _2399_ sky130_fd_sc_hd__a21oi_1
X_3812_ net506 _1640_ VSS VSS VCC VCC _1641_ sky130_fd_sc_hd__and2b_1
X_4792_ _1932_ _2335_ net467 VSS VSS VCC VCC _2336_ sky130_fd_sc_hd__o21ai_1
X_3743_ net700 net76 net390 VSS VSS VCC VCC _0012_ sky130_fd_sc_hd__mux2_1
X_3674_ net530 _1545_ _1546_ _1554_ VSS VSS VCC VCC _1555_ sky130_fd_sc_hd__a31o_2
X_2625_ _0596_ _0597_ _0598_ VSS VSS VCC VCC _0600_ sky130_fd_sc_hd__a21o_1
X_5344_ clknet_4_0__leaf_i_clk _0372_ VSS VSS VCC VCC u_muldiv.divisor\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_2556_ _0525_ _0530_ VSS VSS VCC VCC _0531_ sky130_fd_sc_hd__nor2_1
Xoutput189 net189 VSS VSS VCC VCC o_add[15] sky130_fd_sc_hd__buf_2
X_5275_ clknet_leaf_142_i_clk _0303_ VSS VSS VCC VCC u_muldiv.quotient_msk\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_2487_ net579 net551 VSS VSS VCC VCC _0462_ sky130_fd_sc_hd__nand2_1
X_4226_ u_muldiv.divisor\[3\] _0441_ VSS VSS VCC VCC _1854_ sky130_fd_sc_hd__nor2_1
X_4157_ net552 net499 net192 VSS VSS VCC VCC _0201_ sky130_fd_sc_hd__o21a_1
X_3108_ _1067_ _1068_ VSS VSS VCC VCC _1069_ sky130_fd_sc_hd__nand2_1
X_4088_ u_bits.i_op2\[20\] _1796_ net384 VSS VSS VCC VCC _1797_ sky130_fd_sc_hd__o21ai_1
X_3039_ u_muldiv.dividend\[27\] net419 net364 u_muldiv.o_div\[27\] net442 vssd1 vssd1
+ vccd1 vccd1 _1003_ sky130_fd_sc_hd__a221o_1
Xfanout350 net351 VSS VSS VCC VCC net350 sky130_fd_sc_hd__buf_4
Xfanout361 _0759_ VSS VSS VCC VCC net361 sky130_fd_sc_hd__clkbuf_8
Xfanout372 net373 VSS VSS VCC VCC net372 sky130_fd_sc_hd__clkbuf_4
Xfanout383 net385 VSS VSS VCC VCC net383 sky130_fd_sc_hd__buf_6
Xfanout394 net395 VSS VSS VCC VCC net394 sky130_fd_sc_hd__clkbuf_4
Xinput14 i_csr_data[17] VSS VSS VCC VCC net14 sky130_fd_sc_hd__clkbuf_2
Xinput25 i_csr_data[27] VSS VSS VCC VCC net25 sky130_fd_sc_hd__clkbuf_4
Xinput36 i_csr_data[8] VSS VSS VCC VCC net36 sky130_fd_sc_hd__clkbuf_1
Xinput47 i_op1[11] VSS VSS VCC VCC net47 sky130_fd_sc_hd__clkbuf_1
Xinput58 i_op1[21] VSS VSS VCC VCC net58 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 i_op1[31] VSS VSS VCC VCC net69 sky130_fd_sc_hd__clkbuf_1
X_3390_ _1211_ net522 _0576_ net537 VSS VSS VCC VCC _1288_ sky130_fd_sc_hd__a31o_1
X_5060_ clknet_leaf_58_i_clk _0093_ VSS VSS VCC VCC net244 sky130_fd_sc_hd__dfxtp_2
X_4011_ net602 _1734_ _1735_ VSS VSS VCC VCC _1736_ sky130_fd_sc_hd__a21oi_1
X_4913_ u_muldiv.divisor\[20\] net481 net334 u_muldiv.divisor\[21\] vssd1 vssd1 vccd1
+ vccd1 _0365_ sky130_fd_sc_hd__a22o_1
X_4844_ u_muldiv.dividend\[27\] u_muldiv.dividend\[26\] u_muldiv.dividend\[25\] _2345_
+ VSS VSS VCC VCC _2384_ sky130_fd_sc_hd__or4_1
X_4775_ u_muldiv.dividend\[21\] u_muldiv.dividend\[20\] u_muldiv.dividend\[19\] vssd1
+ vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__nor3_1
X_3726_ net605 _1602_ _1601_ VSS VSS VCC VCC _1603_ sky130_fd_sc_hd__o21a_1
X_3657_ u_bits.i_op2\[16\] net685 net351 _1538_ VSS VSS VCC VCC _1539_ sky130_fd_sc_hd__o211a_1
X_2608_ _0547_ _0559_ _0580_ VSS VSS VCC VCC _0583_ sky130_fd_sc_hd__a21boi_4
X_3588_ net441 u_muldiv.mul\[43\] _0758_ _1474_ VSS VSS VCC VCC _1475_ sky130_fd_sc_hd__a31o_1
X_2539_ _0511_ _0512_ net430 VSS VSS VCC VCC _0514_ sky130_fd_sc_hd__o21ai_1
X_5327_ clknet_leaf_125_i_clk _0355_ VSS VSS VCC VCC u_muldiv.divisor\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_5258_ clknet_leaf_95_i_clk _0286_ VSS VSS VCC VCC u_muldiv.quotient_msk\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4209_ op_cnt\[3\] _1838_ _1839_ VSS VSS VCC VCC _0249_ sky130_fd_sc_hd__o21ba_1
X_5189_ clknet_leaf_97_i_clk _0221_ VSS VSS VCC VCC u_muldiv.mul\[6\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_1_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_2890_ net564 u_bits.i_op2\[23\] net669 VSS VSS VCC VCC _0862_ sky130_fd_sc_hd__nand3b_1
X_4560_ net459 _2123_ _2124_ net498 VSS VSS VCC VCC _2125_ sky130_fd_sc_hd__a31oi_1
X_3511_ net352 _1398_ _1399_ _1401_ net521 VSS VSS VCC VCC _1403_ sky130_fd_sc_hd__a41o_1
X_4491_ net315 _2092_ u_muldiv.o_div\[27\] VSS VSS VCC VCC _2093_ sky130_fd_sc_hd__a21o_1
X_3442_ net678 net676 net674 net671 net641 net634 VSS VSS VCC VCC _1337_ sky130_fd_sc_hd__mux4_1
X_3373_ net675 net672 net671 net668 net638 net631 VSS VSS VCC VCC _1271_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_177_i_clk clknet_4_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_177_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5112_ clknet_leaf_35_i_clk _0145_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_5043_ clknet_leaf_167_i_clk _0076_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_100_i_clk clknet_4_14__leaf_i_clk VSS VSS VCC VCC clknet_leaf_100_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_115_i_clk clknet_4_11__leaf_i_clk VSS VSS VCC VCC clknet_leaf_115_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4827_ net667 net664 net662 _2338_ VSS VSS VCC VCC _2368_ sky130_fd_sc_hd__or4_1
X_4758_ u_muldiv.dividend\[20\] u_muldiv.dividend\[19\] _0450_ _2280_ vssd1 vssd1
+ vccd1 vccd1 _2305_ sky130_fd_sc_hd__and4bb_1
X_3709_ net604 _1365_ net327 VSS VSS VCC VCC _1587_ sky130_fd_sc_hd__o21a_1
X_4689_ u_muldiv.dividend\[14\] u_muldiv.dividend\[13\] _2222_ VSS VSS VCC VCC
+ _2242_ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_94_i_clk clknet_4_14__leaf_i_clk VSS VSS VCC VCC clknet_leaf_94_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_32_i_clk clknet_4_4__leaf_i_clk VSS VSS VCC VCC clknet_leaf_32_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3991_ net433 net465 VSS VSS VCC VCC _1720_ sky130_fd_sc_hd__nand2_8
X_2942_ net611 _0903_ _0911_ VSS VSS VCC VCC _0912_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_47_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_47_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2873_ net704 net707 net708 net711 net644 net635 VSS VSS VCC VCC _0845_ sky130_fd_sc_hd__mux4_1
X_4612_ net710 net708 net706 _2143_ VSS VSS VCC VCC _2172_ sky130_fd_sc_hd__or4b_2
X_4543_ u_muldiv.dividend\[0\] net464 VSS VSS VCC VCC _2109_ sky130_fd_sc_hd__xnor2_1
X_4474_ net317 _2079_ u_muldiv.o_div\[23\] VSS VSS VCC VCC _2080_ sky130_fd_sc_hd__a21oi_1
X_3425_ _1320_ net606 VSS VSS VCC VCC _1321_ sky130_fd_sc_hd__nand2b_1
X_3356_ net568 u_wr_mux.i_reg_data2\[28\] net416 net305 VSS VSS VCC VCC _1262_
+ sky130_fd_sc_hd__a22o_2
X_3287_ _1205_ _1218_ VSS VSS VCC VCC _1219_ sky130_fd_sc_hd__nand2_2
X_5026_ clknet_leaf_49_i_clk _0059_ VSS VSS VCC VCC u_bits.i_op2\[15\] sky130_fd_sc_hd__dfxtp_4
X_3210_ _0544_ _0546_ _0560_ _0579_ _0580_ VSS VSS VCC VCC _1162_ sky130_fd_sc_hd__o2111ai_4
X_4190_ u_muldiv.mul\[20\] u_muldiv.mul\[19\] net404 VSS VSS VCC VCC _0234_
+ sky130_fd_sc_hd__mux2_1
X_3141_ _1029_ _1068_ _1067_ VSS VSS VCC VCC _1100_ sky130_fd_sc_hd__a21bo_1
X_3072_ _1034_ _1033_ VSS VSS VCC VCC _1035_ sky130_fd_sc_hd__nor2_1
X_3974_ u_wr_mux.i_reg_data2\[18\] net153 net386 VSS VSS VCC VCC _0136_ sky130_fd_sc_hd__mux2_1
X_2925_ net601 _0894_ net327 VSS VSS VCC VCC _0895_ sky130_fd_sc_hd__o21ai_1
X_2856_ _0825_ _0826_ _0822_ VSS VSS VCC VCC _0829_ sky130_fd_sc_hd__a21o_1
X_2787_ u_muldiv.mul\[54\] net363 net357 u_muldiv.mul\[22\] _0756_ vssd1 vssd1 vccd1
+ vccd1 _0761_ sky130_fd_sc_hd__a221o_2
X_4526_ u_muldiv.quotient_msk\[14\] net491 net338 u_muldiv.quotient_msk\[15\] vssd1
+ vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__a22o_1
X_4457_ u_muldiv.o_div\[18\] u_muldiv.o_div\[19\] u_muldiv.o_div\[20\] _2058_ vssd1
+ vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__or4_2
Xfanout702 net703 VSS VSS VCC VCC net702 sky130_fd_sc_hd__buf_2
Xfanout713 net714 VSS VSS VCC VCC net713 sky130_fd_sc_hd__buf_4
X_3408_ net565 net717 net632 VSS VSS VCC VCC _1305_ sky130_fd_sc_hd__nand3b_1
Xfanout724 _1608_ VSS VSS VCC VCC net724 sky130_fd_sc_hd__clkbuf_4
Xfanout735 net38 VSS VSS VCC VCC net735 sky130_fd_sc_hd__buf_12
X_4388_ net320 _2009_ _2011_ VSS VSS VCC VCC _0256_ sky130_fd_sc_hd__a21oi_1
X_3339_ u_wr_mux.i_reg_data2\[15\] net308 net417 VSS VSS VCC VCC net285 sky130_fd_sc_hd__mux2_8
X_5009_ clknet_leaf_24_i_clk _0042_ VSS VSS VCC VCC u_pc_sel.i_inst_jal_jalr
+ sky130_fd_sc_hd__dfxtp_2
X_2710_ _0662_ _0684_ VSS VSS VCC VCC _0685_ sky130_fd_sc_hd__nor2_1
X_3690_ net731 net15 _1569_ VSS VSS VCC VCC net254 sky130_fd_sc_hd__o21a_4
X_2641_ net648 net554 net707 net539 net425 VSS VSS VCC VCC _0616_ sky130_fd_sc_hd__o2111ai_4
Xoutput305 net305 VSS VSS VCC VCC o_wdata[4] sky130_fd_sc_hd__buf_2
X_2572_ net431 _0541_ _0546_ VSS VSS VCC VCC _0547_ sky130_fd_sc_hd__a21o_1
X_5360_ clknet_leaf_102_i_clk _0387_ VSS VSS VCC VCC u_muldiv.mul\[39\] sky130_fd_sc_hd__dfxtp_1
X_4311_ u_muldiv.divisor\[21\] u_muldiv.dividend\[21\] VSS VSS VCC VCC _1939_
+ sky130_fd_sc_hd__and2b_1
X_5291_ clknet_leaf_112_i_clk _0319_ VSS VSS VCC VCC u_muldiv.dividend\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_4242_ u_muldiv.divisor\[6\] _0443_ _1845_ VSS VSS VCC VCC _1870_ sky130_fd_sc_hd__or3b_1
X_4173_ u_muldiv.mul\[3\] u_muldiv.mul\[2\] net404 VSS VSS VCC VCC _0217_
+ sky130_fd_sc_hd__mux2_1
X_3124_ net560 _1083_ VSS VSS VCC VCC _1084_ sky130_fd_sc_hd__or2_1
X_3055_ net659 net582 net411 _1018_ VSS VSS VCC VCC _1019_ sky130_fd_sc_hd__a31o_1
X_3957_ net290 net155 net392 VSS VSS VCC VCC _0119_ sky130_fd_sc_hd__mux2_1
X_2908_ _0749_ _0878_ VSS VSS VCC VCC _0879_ sky130_fd_sc_hd__nor2_2
X_3888_ net501 _1697_ VSS VSS VCC VCC _1698_ sky130_fd_sc_hd__and2b_1
X_2839_ net453 _0812_ _0807_ _0811_ VSS VSS VCC VCC _0813_ sky130_fd_sc_hd__a211o_1
X_4509_ u_muldiv.quotient_msk\[31\] net434 _2103_ VSS VSS VCC VCC _2107_ sky130_fd_sc_hd__a21o_1
Xfanout510 net511 VSS VSS VCC VCC net510 sky130_fd_sc_hd__clkbuf_2
Xfanout521 net522 VSS VSS VCC VCC net521 sky130_fd_sc_hd__buf_6
Xfanout532 net543 VSS VSS VCC VCC net532 sky130_fd_sc_hd__buf_4
Xfanout543 net544 VSS VSS VCC VCC net543 sky130_fd_sc_hd__clkbuf_8
Xfanout554 net555 VSS VSS VCC VCC net554 sky130_fd_sc_hd__clkbuf_16
Xfanout565 net568 VSS VSS VCC VCC net565 sky130_fd_sc_hd__clkbuf_4
Xfanout576 net243 VSS VSS VCC VCC net576 sky130_fd_sc_hd__clkbuf_8
Xfanout587 u_bits.i_op2\[19\] VSS VSS VCC VCC net587 sky130_fd_sc_hd__buf_8
Xfanout598 u_bits.i_op2\[7\] VSS VSS VCC VCC net598 sky130_fd_sc_hd__buf_6
X_4860_ _1966_ _1960_ _1964_ VSS VSS VCC VCC _2398_ sky130_fd_sc_hd__o21bai_1
X_3811_ net597 net599 net545 VSS VSS VCC VCC _1640_ sky130_fd_sc_hd__mux2_1
X_4791_ _1928_ _2326_ _1926_ VSS VSS VCC VCC _2335_ sky130_fd_sc_hd__a21oi_1
X_3742_ net703 net75 net396 VSS VSS VCC VCC _0011_ sky130_fd_sc_hd__mux2_1
X_3673_ net356 _1221_ _1553_ net520 net444 VSS VSS VCC VCC _1554_ sky130_fd_sc_hd__o221a_1
X_2624_ _0596_ _0597_ _0598_ VSS VSS VCC VCC _0599_ sky130_fd_sc_hd__a21oi_1
X_5343_ clknet_leaf_173_i_clk _0371_ VSS VSS VCC VCC u_muldiv.divisor\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_2555_ _0524_ _0523_ _0522_ VSS VSS VCC VCC _0530_ sky130_fd_sc_hd__and3b_2
X_5274_ clknet_leaf_139_i_clk _0302_ VSS VSS VCC VCC u_muldiv.quotient_msk\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_2486_ net579 net551 VSS VSS VCC VCC _0461_ sky130_fd_sc_hd__nand2b_1
X_4225_ _0441_ u_muldiv.divisor\[3\] VSS VSS VCC VCC _1853_ sky130_fd_sc_hd__nand2_1
X_4156_ net552 net500 net191 VSS VSS VCC VCC _0200_ sky130_fd_sc_hd__o21a_1
X_3107_ _1065_ _1066_ _1063_ _1064_ VSS VSS VCC VCC _1068_ sky130_fd_sc_hd__o211ai_2
X_4087_ u_bits.i_op2\[18\] net587 _1787_ net380 VSS VSS VCC VCC _1796_ sky130_fd_sc_hd__o31a_1
X_3038_ _1002_ VSS VSS VCC VCC net202 sky130_fd_sc_hd__clkinv_4
X_4989_ clknet_leaf_34_i_clk _0022_ VSS VSS VCC VCC u_bits.i_op1\[19\] sky130_fd_sc_hd__dfxtp_4
Xfanout340 net341 VSS VSS VCC VCC net340 sky130_fd_sc_hd__buf_2
Xfanout351 _0785_ VSS VSS VCC VCC net351 sky130_fd_sc_hd__buf_4
Xfanout362 net363 VSS VSS VCC VCC net362 sky130_fd_sc_hd__clkbuf_2
Xfanout373 net374 VSS VSS VCC VCC net373 sky130_fd_sc_hd__clkbuf_4
Xfanout384 net385 VSS VSS VCC VCC net384 sky130_fd_sc_hd__buf_4
Xfanout395 _1610_ VSS VSS VCC VCC net395 sky130_fd_sc_hd__buf_6
Xinput15 i_csr_data[18] VSS VSS VCC VCC net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 i_csr_data[28] VSS VSS VCC VCC net26 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput37 i_csr_data[9] VSS VSS VCC VCC net37 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput48 i_op1[12] VSS VSS VCC VCC net48 sky130_fd_sc_hd__clkbuf_1
Xinput59 i_op1[22] VSS VSS VCC VCC net59 sky130_fd_sc_hd__clkbuf_1
X_4010_ net602 _1734_ net383 VSS VSS VCC VCC _1735_ sky130_fd_sc_hd__o21ai_1
X_4912_ u_muldiv.divisor\[19\] net481 net334 u_muldiv.divisor\[20\] vssd1 vssd1 vccd1
+ vccd1 _0364_ sky130_fd_sc_hd__a22o_1
X_4843_ net433 _2381_ _2382_ net332 VSS VSS VCC VCC _2383_ sky130_fd_sc_hd__a31oi_2
X_4774_ _2314_ _2315_ net467 _2319_ VSS VSS VCC VCC _2320_ sky130_fd_sc_hd__a31oi_1
X_3725_ _0938_ _0942_ _0944_ _0947_ net454 net451 VSS VSS VCC VCC _1602_ sky130_fd_sc_hd__mux4_1
X_3656_ _0428_ net564 net685 VSS VSS VCC VCC _1538_ sky130_fd_sc_hd__or3b_1
X_2607_ _0568_ _0578_ _0581_ _0562_ VSS VSS VCC VCC _0582_ sky130_fd_sc_hd__nand4_4
X_3587_ u_muldiv.dividend\[11\] net420 net368 u_muldiv.o_div\[11\] net360 vssd1 vssd1
+ vccd1 vccd1 _1474_ sky130_fd_sc_hd__a221o_2
X_5326_ clknet_leaf_125_i_clk _0354_ VSS VSS VCC VCC u_muldiv.divisor\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2538_ net535 net683 _0463_ _0511_ net427 VSS VSS VCC VCC _0513_ sky130_fd_sc_hd__a311oi_1
X_5257_ clknet_leaf_95_i_clk _0285_ VSS VSS VCC VCC u_muldiv.quotient_msk\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2469_ u_muldiv.dividend\[4\] VSS VSS VCC VCC _0444_ sky130_fd_sc_hd__clkinv_2
X_4208_ op_cnt\[0\] op_cnt\[1\] op_cnt\[2\] op_cnt\[3\] net510 VSS VSS VCC VCC
+ _1839_ sky130_fd_sc_hd__a41o_1
X_5188_ clknet_leaf_97_i_clk _0220_ VSS VSS VCC VCC u_muldiv.mul\[5\] sky130_fd_sc_hd__dfxtp_1
X_4139_ u_muldiv.quotient_msk\[31\] net477 net383 VSS VSS VCC VCC _0183_ sky130_fd_sc_hd__a21o_1
Xclkbuf_4_12__f_i_clk clknet_2_3_0_i_clk VSS VSS VCC VCC clknet_4_12__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3510_ u_bits.i_op2\[6\] net706 net353 VSS VSS VCC VCC _1402_ sky130_fd_sc_hd__a21oi_1
X_4490_ u_muldiv.quotient_msk\[27\] net433 _2088_ VSS VSS VCC VCC _2092_ sky130_fd_sc_hd__a21o_1
X_3441_ net578 u_pc_sel.i_pc_next\[2\] _1335_ _1336_ VSS VSS VCC VCC net267
+ sky130_fd_sc_hd__a22o_1
X_3372_ net684 net683 net679 net677 net637 net627 VSS VSS VCC VCC _1270_ sky130_fd_sc_hd__mux4_2
X_5111_ clknet_leaf_90_i_clk _0144_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[26\]
+ sky130_fd_sc_hd__dfxtp_2
X_5042_ clknet_leaf_11_i_clk _0075_ VSS VSS VCC VCC u_bits.i_op2\[31\] sky130_fd_sc_hd__dfxtp_4
X_4826_ _2365_ _1957_ _1950_ VSS VSS VCC VCC _2367_ sky130_fd_sc_hd__a21o_1
X_4757_ u_muldiv.dividend\[19\] u_muldiv.dividend\[18\] net462 _2262_ u_muldiv.dividend\[20\]
+ VSS VSS VCC VCC _2304_ sky130_fd_sc_hd__o41a_1
X_3708_ net565 _1585_ net558 net572 VSS VSS VCC VCC _1586_ sky130_fd_sc_hd__or4b_1
X_4688_ u_muldiv.dividend\[13\] _2241_ net321 VSS VSS VCC VCC _0326_ sky130_fd_sc_hd__mux2_1
X_3639_ net608 net452 _0838_ _1521_ _0765_ VSS VSS VCC VCC _1522_ sky130_fd_sc_hd__o311a_1
X_5309_ clknet_leaf_167_i_clk _0337_ VSS VSS VCC VCC u_muldiv.dividend\[24\]
+ sky130_fd_sc_hd__dfxtp_2
X_3990_ net490 net459 VSS VSS VCC VCC _1719_ sky130_fd_sc_hd__nor2_1
X_2941_ net346 _0906_ _0905_ _0904_ net345 VSS VSS VCC VCC _0911_ sky130_fd_sc_hd__o221a_1
X_2872_ net609 _0843_ net328 VSS VSS VCC VCC _0844_ sky130_fd_sc_hd__o21a_1
X_4611_ net708 net706 VSS VSS VCC VCC _2171_ sky130_fd_sc_hd__nor2_1
X_4542_ u_muldiv.quotient_msk\[30\] net477 net333 u_muldiv.quotient_msk\[31\] vssd1
+ vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__a22o_1
X_4473_ _2074_ u_muldiv.quotient_msk\[23\] net434 VSS VSS VCC VCC _2079_ sky130_fd_sc_hd__mux2_1
X_3424_ _0770_ _0776_ _1319_ _0771_ net615 net456 VSS VSS VCC VCC _1320_ sky130_fd_sc_hd__mux4_2
X_3355_ u_wr_mux.i_reg_data2\[11\] _0764_ _1261_ VSS VSS VCC VCC net298 sky130_fd_sc_hd__a21o_4
X_3286_ _0525_ _0530_ _0741_ _0732_ VSS VSS VCC VCC _1218_ sky130_fd_sc_hd__o211ai_2
X_5025_ clknet_leaf_26_i_clk _0058_ VSS VSS VCC VCC u_bits.i_op2\[14\] sky130_fd_sc_hd__dfxtp_4
X_4809_ net466 _2350_ _2351_ _2348_ _2347_ VSS VSS VCC VCC _2352_ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_161_i_clk clknet_4_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_161_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_114_i_clk clknet_4_11__leaf_i_clk VSS VSS VCC VCC clknet_leaf_114_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3140_ _1034_ _1033_ _1097_ VSS VSS VCC VCC _1099_ sky130_fd_sc_hd__o21bai_1
X_3071_ _0998_ _0966_ _0968_ _1031_ _0996_ VSS VSS VCC VCC _1034_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_129_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_129_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3973_ u_wr_mux.i_reg_data2\[17\] net152 net391 VSS VSS VCC VCC _0135_ sky130_fd_sc_hd__mux2_1
X_2924_ net611 _0893_ net347 VSS VSS VCC VCC _0894_ sky130_fd_sc_hd__o21a_1
X_2855_ _0822_ _0825_ _0826_ VSS VSS VCC VCC _0828_ sky130_fd_sc_hd__nand3_1
X_2786_ net559 net414 VSS VSS VCC VCC _0760_ sky130_fd_sc_hd__nor2_8
X_4525_ u_muldiv.quotient_msk\[13\] net491 net340 u_muldiv.quotient_msk\[14\] vssd1
+ vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__a22o_1
X_4456_ net322 _2063_ _2065_ u_muldiv.o_div\[19\] VSS VSS VCC VCC _0270_ sky130_fd_sc_hd__o22a_1
Xfanout703 u_bits.i_op1\[8\] VSS VSS VCC VCC net703 sky130_fd_sc_hd__buf_6
X_3407_ _0907_ net345 _0936_ VSS VSS VCC VCC _1304_ sky130_fd_sc_hd__and3_1
Xfanout714 u_bits.i_op1\[3\] VSS VSS VCC VCC net714 sky130_fd_sc_hd__buf_4
X_4387_ net320 _2010_ u_muldiv.o_div\[5\] VSS VSS VCC VCC _2011_ sky130_fd_sc_hd__a21oi_1
Xfanout725 net726 VSS VSS VCC VCC net725 sky130_fd_sc_hd__clkbuf_4
X_3338_ u_wr_mux.i_reg_data2\[14\] net307 net418 VSS VSS VCC VCC net284 sky130_fd_sc_hd__mux2_4
X_3269_ _1206_ _0509_ _0506_ VSS VSS VCC VCC _1207_ sky130_fd_sc_hd__a21boi_2
X_5008_ clknet_leaf_30_i_clk _0041_ VSS VSS VCC VCC net239 sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_93_i_clk clknet_4_14__leaf_i_clk VSS VSS VCC VCC clknet_leaf_93_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_31_i_clk clknet_4_4__leaf_i_clk VSS VSS VCC VCC clknet_leaf_31_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_4_0__f_i_clk clknet_2_0_0_i_clk VSS VSS VCC VCC clknet_4_0__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_46_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_46_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2640_ _0613_ _0612_ _0611_ VSS VSS VCC VCC _0615_ sky130_fd_sc_hd__nand3b_4
X_2571_ _0545_ _0536_ VSS VSS VCC VCC _0546_ sky130_fd_sc_hd__nand2_2
Xoutput306 net306 VSS VSS VCC VCC o_wdata[5] sky130_fd_sc_hd__buf_2
X_4310_ u_muldiv.dividend\[21\] u_muldiv.divisor\[21\] VSS VSS VCC VCC _1938_
+ sky130_fd_sc_hd__nand2b_1
X_5290_ clknet_leaf_96_i_clk _0318_ VSS VSS VCC VCC u_muldiv.dividend\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_4241_ u_muldiv.divisor\[6\] _0443_ _1868_ VSS VSS VCC VCC _1869_ sky130_fd_sc_hd__o21a_1
X_4172_ u_muldiv.mul\[2\] u_muldiv.mul\[1\] net404 VSS VSS VCC VCC _0216_
+ sky130_fd_sc_hd__mux2_1
X_3123_ net655 net581 VSS VSS VCC VCC _1083_ sky130_fd_sc_hd__nand2_1
X_3054_ net659 net582 _1017_ net348 VSS VSS VCC VCC _1018_ sky130_fd_sc_hd__o211a_1
X_3956_ net279 net144 net395 VSS VSS VCC VCC _0118_ sky130_fd_sc_hd__mux2_1
X_2907_ _0470_ _0472_ _0828_ _0829_ VSS VSS VCC VCC _0878_ sky130_fd_sc_hd__nand4_1
X_3887_ net582 net584 net545 VSS VSS VCC VCC _1697_ sky130_fd_sc_hd__mux2_1
X_2838_ net670 net673 net675 net677 net638 net627 VSS VSS VCC VCC _0812_ sky130_fd_sc_hd__mux4_2
X_2769_ _0732_ _0741_ VSS VSS VCC VCC _0744_ sky130_fd_sc_hd__nand2_4
X_4508_ u_muldiv.o_div\[31\] _2103_ net477 net466 VSS VSS VCC VCC _2106_ sky130_fd_sc_hd__o2bb2a_1
X_4439_ u_muldiv.o_div\[16\] _2050_ _2051_ VSS VSS VCC VCC _2052_ sky130_fd_sc_hd__a21boi_1
Xfanout500 u_muldiv.i_on_wait VSS VSS VCC VCC net500 sky130_fd_sc_hd__buf_6
Xfanout511 net240 VSS VSS VCC VCC net511 sky130_fd_sc_hd__buf_2
Xfanout522 u_mux.i_add_override VSS VSS VCC VCC net522 sky130_fd_sc_hd__buf_6
Xfanout533 net536 VSS VSS VCC VCC net533 sky130_fd_sc_hd__clkbuf_4
Xfanout544 u_mux.i_group_mux VSS VSS VCC VCC net544 sky130_fd_sc_hd__buf_8
Xfanout555 u_muldiv.i_is_div VSS VSS VCC VCC net555 sky130_fd_sc_hd__buf_8
Xfanout566 net567 VSS VSS VCC VCC net566 sky130_fd_sc_hd__clkbuf_4
Xfanout577 net578 VSS VSS VCC VCC net577 sky130_fd_sc_hd__clkbuf_8
Xfanout588 u_bits.i_op2\[18\] VSS VSS VCC VCC net588 sky130_fd_sc_hd__buf_6
Xfanout599 u_bits.i_op2\[6\] VSS VSS VCC VCC net599 sky130_fd_sc_hd__clkbuf_4
X_3810_ net599 net725 _1639_ _1638_ VSS VSS VCC VCC _0050_ sky130_fd_sc_hd__o22a_1
X_4790_ u_muldiv.dividend\[22\] _2334_ net317 VSS VSS VCC VCC _0335_ sky130_fd_sc_hd__mux2_1
X_3741_ u_bits.i_op1\[7\] net74 net389 VSS VSS VCC VCC _0010_ sky130_fd_sc_hd__mux2_1
X_3672_ net409 _1549_ _1552_ _1547_ VSS VSS VCC VCC _1553_ sky130_fd_sc_hd__o211a_1
X_2623_ net709 u_muldiv.add_prev\[5\] net539 VSS VSS VCC VCC _0598_ sky130_fd_sc_hd__mux2_2
X_5342_ clknet_leaf_172_i_clk _0370_ VSS VSS VCC VCC u_muldiv.divisor\[25\]
+ sky130_fd_sc_hd__dfxtp_2
X_2554_ _0518_ _0519_ VSS VSS VCC VCC _0529_ sky130_fd_sc_hd__nand2_2
X_5273_ clknet_4_10__leaf_i_clk _0301_ VSS VSS VCC VCC u_muldiv.quotient_msk\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_2485_ net579 net551 VSS VSS VCC VCC _0460_ sky130_fd_sc_hd__and2b_2
X_4224_ _0441_ u_muldiv.divisor\[3\] VSS VSS VCC VCC _1852_ sky130_fd_sc_hd__and2_1
X_4155_ _1205_ _1218_ net401 VSS VSS VCC VCC _0199_ sky130_fd_sc_hd__and3_1
X_3106_ net533 u_muldiv.add_prev\[29\] _1063_ _1064_ _1066_ VSS VSS VCC VCC
+ _1067_ sky130_fd_sc_hd__a221o_1
X_4086_ net590 _1794_ net589 _1780_ VSS VSS VCC VCC _1795_ sky130_fd_sc_hd__or4_1
X_3037_ _1000_ _1001_ VSS VSS VCC VCC _1002_ sky130_fd_sc_hd__nand2_1
X_4988_ clknet_leaf_0_i_clk _0021_ VSS VSS VCC VCC u_bits.i_op1\[18\] sky130_fd_sc_hd__dfxtp_1
X_3939_ net234 net138 net393 VSS VSS VCC VCC _0102_ sky130_fd_sc_hd__mux2_1
Xfanout330 net331 VSS VSS VCC VCC net330 sky130_fd_sc_hd__buf_6
Xfanout341 net344 VSS VSS VCC VCC net341 sky130_fd_sc_hd__buf_4
Xfanout352 _0783_ VSS VSS VCC VCC net352 sky130_fd_sc_hd__buf_4
Xfanout363 _0759_ VSS VSS VCC VCC net363 sky130_fd_sc_hd__buf_6
Xfanout374 _2113_ VSS VSS VCC VCC net374 sky130_fd_sc_hd__buf_6
Xfanout385 _1721_ VSS VSS VCC VCC net385 sky130_fd_sc_hd__clkbuf_16
Xfanout396 net397 VSS VSS VCC VCC net396 sky130_fd_sc_hd__buf_4
Xinput16 i_csr_data[19] VSS VSS VCC VCC net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 i_csr_data[29] VSS VSS VCC VCC net27 sky130_fd_sc_hd__clkbuf_2
Xinput38 i_csr_read VSS VSS VCC VCC net38 sky130_fd_sc_hd__buf_4
Xinput49 i_op1[13] VSS VSS VCC VCC net49 sky130_fd_sc_hd__clkbuf_1
X_4911_ u_muldiv.divisor\[18\] net488 net341 u_muldiv.divisor\[19\] vssd1 vssd1 vccd1
+ vccd1 _0363_ sky130_fd_sc_hd__a22o_1
X_4842_ _2380_ net369 net658 VSS VSS VCC VCC _2382_ sky130_fd_sc_hd__a21o_1
X_4773_ net481 _2317_ _2318_ _1720_ VSS VSS VCC VCC _2319_ sky130_fd_sc_hd__o31a_1
X_3724_ net614 _1081_ net604 VSS VSS VCC VCC _1601_ sky130_fd_sc_hd__o21ai_1
X_3655_ _0806_ _0903_ _1536_ VSS VSS VCC VCC _1537_ sky130_fd_sc_hd__a21oi_2
X_2606_ _0544_ _0546_ _0580_ VSS VSS VCC VCC _0581_ sky130_fd_sc_hd__o21a_1
X_3586_ net521 _1472_ _0762_ _1188_ VSS VSS VCC VCC _1473_ sky130_fd_sc_hd__o22a_1
X_5325_ clknet_4_10__leaf_i_clk _0353_ VSS VSS VCC VCC u_muldiv.divisor\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_2537_ _0459_ net423 net535 net683 VSS VSS VCC VCC _0512_ sky130_fd_sc_hd__and4_1
X_5256_ clknet_leaf_94_i_clk _0284_ VSS VSS VCC VCC u_muldiv.quotient_msk\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2468_ u_muldiv.dividend\[6\] VSS VSS VCC VCC _0443_ sky130_fd_sc_hd__clkinv_2
X_4207_ net510 _1837_ _1838_ VSS VSS VCC VCC _0248_ sky130_fd_sc_hd__nor3_1
X_5187_ clknet_leaf_97_i_clk _0219_ VSS VSS VCC VCC u_muldiv.mul\[4\] sky130_fd_sc_hd__dfxtp_1
X_4138_ _1835_ net383 net579 net478 u_muldiv.divisor\[62\] VSS VSS VCC VCC
+ _0182_ sky130_fd_sc_hd__a32o_1
X_4069_ _1780_ net380 net590 net329 VSS VSS VCC VCC _1782_ sky130_fd_sc_hd__a31o_1
X_3440_ net28 net731 net578 VSS VSS VCC VCC _1336_ sky130_fd_sc_hd__o21ba_1
X_3371_ net440 _1268_ VSS VSS VCC VCC _1269_ sky130_fd_sc_hd__nand2_2
X_5110_ clknet_leaf_84_i_clk _0143_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[25\]
+ sky130_fd_sc_hd__dfxtp_4
X_5041_ clknet_leaf_56_i_clk _0074_ VSS VSS VCC VCC u_bits.i_op2\[30\] sky130_fd_sc_hd__dfxtp_1
X_4825_ _1950_ _2365_ _1957_ VSS VSS VCC VCC _2366_ sky130_fd_sc_hd__nand3_1
X_4756_ u_muldiv.dividend\[19\] _1993_ _2303_ VSS VSS VCC VCC _0332_ sky130_fd_sc_hd__o21a_1
X_3707_ net613 _1045_ _1049_ _0806_ _1584_ VSS VSS VCC VCC _1585_ sky130_fd_sc_hd__a221o_1
X_4687_ _2239_ _2240_ _2238_ VSS VSS VCC VCC _2241_ sky130_fd_sc_hd__a21o_1
X_3638_ _0842_ net347 net608 VSS VSS VCC VCC _1521_ sky130_fd_sc_hd__a21bo_1
X_3569_ u_bits.i_op2\[10\] net697 net352 VSS VSS VCC VCC _1457_ sky130_fd_sc_hd__a21oi_1
X_5308_ clknet_4_2__leaf_i_clk _0336_ VSS VSS VCC VCC u_muldiv.dividend\[23\]
+ sky130_fd_sc_hd__dfxtp_2
X_5239_ clknet_leaf_130_i_clk _0267_ VSS VSS VCC VCC u_muldiv.o_div\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_2940_ net610 net565 net558 net572 VSS VSS VCC VCC _0910_ sky130_fd_sc_hd__or4b_4
X_2871_ _0838_ _0842_ net616 VSS VSS VCC VCC _0843_ sky130_fd_sc_hd__mux2_1
X_4610_ _1869_ _1872_ net470 VSS VSS VCC VCC _2170_ sky130_fd_sc_hd__o21ai_1
X_4541_ u_muldiv.quotient_msk\[29\] net477 net334 u_muldiv.quotient_msk\[30\] vssd1
+ vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__a22o_1
X_4472_ _2074_ net480 u_muldiv.o_div\[23\] net383 VSS VSS VCC VCC _2078_ sky130_fd_sc_hd__a31o_1
X_3423_ net680 net677 net676 net674 net639 net632 VSS VSS VCC VCC _1319_ sky130_fd_sc_hd__mux4_1
X_3354_ net563 u_wr_mux.i_reg_data2\[27\] net416 net304 VSS VSS VCC VCC _1261_
+ sky130_fd_sc_hd__a22o_1
X_3285_ _1175_ _1216_ _1183_ _1177_ VSS VSS VCC VCC _1217_ sky130_fd_sc_hd__nand4_1
X_5024_ clknet_leaf_14_i_clk _0057_ VSS VSS VCC VCC u_bits.i_op2\[13\] sky130_fd_sc_hd__dfxtp_4
X_4808_ net667 _2338_ net369 net664 VSS VSS VCC VCC _2351_ sky130_fd_sc_hd__o211a_1
X_4739_ _2286_ net469 VSS VSS VCC VCC _2288_ sky130_fd_sc_hd__nand2_1
X_3070_ _0882_ _0885_ _1032_ VSS VSS VCC VCC _1033_ sky130_fd_sc_hd__a21oi_2
X_3972_ u_wr_mux.i_reg_data2\[16\] net151 net393 VSS VSS VCC VCC _0134_ sky130_fd_sc_hd__mux2_1
X_2923_ _0891_ _0892_ net624 VSS VSS VCC VCC _0893_ sky130_fd_sc_hd__mux2_1
X_2854_ _0822_ _0825_ _0826_ VSS VSS VCC VCC _0827_ sky130_fd_sc_hd__and3_1
X_2785_ net560 net570 net440 VSS VSS VCC VCC _0759_ sky130_fd_sc_hd__o21a_4
X_4524_ u_muldiv.quotient_msk\[12\] net492 net339 u_muldiv.quotient_msk\[13\] vssd1
+ vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__a22o_1
X_4455_ net324 net375 _2060_ _2064_ VSS VSS VCC VCC _2065_ sky130_fd_sc_hd__o2bb2a_1
X_3406_ _1302_ _1299_ _1295_ _0933_ net611 net605 VSS VSS VCC VCC _1303_ sky130_fd_sc_hd__mux4_1
Xfanout704 net705 VSS VSS VCC VCC net704 sky130_fd_sc_hd__buf_4
X_4386_ _2006_ u_muldiv.quotient_msk\[5\] net438 VSS VSS VCC VCC _2010_ sky130_fd_sc_hd__mux2_1
Xfanout715 u_bits.i_op1\[2\] VSS VSS VCC VCC net715 sky130_fd_sc_hd__buf_4
Xfanout726 _1608_ VSS VSS VCC VCC net726 sky130_fd_sc_hd__buf_2
X_3337_ u_wr_mux.i_reg_data2\[13\] net306 net416 VSS VSS VCC VCC net283 sky130_fd_sc_hd__mux2_8
X_3268_ _0744_ _0532_ _0526_ VSS VSS VCC VCC _1206_ sky130_fd_sc_hd__a21bo_2
X_5007_ clknet_leaf_46_i_clk _0040_ VSS VSS VCC VCC net238 sky130_fd_sc_hd__dfxtp_4
X_3199_ _1142_ _1154_ net735 VSS VSS VCC VCC _1155_ sky130_fd_sc_hd__a21oi_4
X_2570_ _0421_ net538 net518 net525 _0540_ VSS VSS VCC VCC _0545_ sky130_fd_sc_hd__o221ai_2
Xoutput307 net307 VSS VSS VCC VCC o_wdata[6] sky130_fd_sc_hd__buf_2
X_4240_ _1866_ _1867_ VSS VSS VCC VCC _1868_ sky130_fd_sc_hd__nand2b_1
X_4171_ u_muldiv.mul\[1\] u_muldiv.mul\[0\] net403 VSS VSS VCC VCC _0215_
+ sky130_fd_sc_hd__mux2_1
X_3122_ _0936_ _0937_ _0938_ _0942_ net454 net451 VSS VSS VCC VCC _1082_ sky130_fd_sc_hd__mux4_2
X_3053_ net561 net582 net659 VSS VSS VCC VCC _1017_ sky130_fd_sc_hd__nand3b_1
X_3955_ net278 net507 net726 _1717_ VSS VSS VCC VCC _0117_ sky130_fd_sc_hd__o211a_1
X_2906_ _0876_ VSS VSS VCC VCC _0877_ sky130_fd_sc_hd__inv_2
X_3886_ net584 net725 _1696_ _1695_ VSS VSS VCC VCC _0069_ sky130_fd_sc_hd__o22a_1
X_2837_ _0810_ net619 VSS VSS VCC VCC _0811_ sky130_fd_sc_hd__and2_1
X_2768_ _0638_ _0729_ _0742_ VSS VSS VCC VCC _0743_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_leaf_160_i_clk clknet_4_2__leaf_i_clk VSS VSS VCC VCC clknet_leaf_160_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4507_ u_muldiv.o_div\[30\] net316 _2105_ VSS VSS VCC VCC _0281_ sky130_fd_sc_hd__o21a_1
X_2699_ _0672_ _0673_ net428 VSS VSS VCC VCC _0674_ sky130_fd_sc_hd__a21oi_2
X_4438_ u_muldiv.o_div\[16\] _2050_ net491 VSS VSS VCC VCC _2051_ sky130_fd_sc_hd__o21a_1
Xfanout501 net503 VSS VSS VCC VCC net501 sky130_fd_sc_hd__buf_2
Xfanout512 net513 VSS VSS VCC VCC net512 sky130_fd_sc_hd__buf_2
Xfanout523 alu_ctrl\[2\] VSS VSS VCC VCC net523 sky130_fd_sc_hd__buf_6
Xfanout534 net536 VSS VSS VCC VCC net534 sky130_fd_sc_hd__clkbuf_2
X_4369_ net496 _1994_ _1995_ _1996_ VSS VSS VCC VCC _1997_ sky130_fd_sc_hd__a31o_1
Xfanout545 net547 VSS VSS VCC VCC net545 sky130_fd_sc_hd__buf_4
Xfanout556 net557 VSS VSS VCC VCC net556 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_175_i_clk clknet_4_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_175_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout567 net568 VSS VSS VCC VCC net567 sky130_fd_sc_hd__clkbuf_2
Xfanout578 net243 VSS VSS VCC VCC net578 sky130_fd_sc_hd__buf_6
Xfanout589 u_bits.i_op2\[17\] VSS VSS VCC VCC net589 sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_128_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_128_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3740_ u_bits.i_op1\[6\] net73 net387 VSS VSS VCC VCC _0009_ sky130_fd_sc_hd__mux2_1
X_3671_ u_bits.i_op2\[17\] net683 _0782_ _1551_ VSS VSS VCC VCC _1552_ sky130_fd_sc_hd__a31oi_4
X_2622_ _0594_ _0595_ net431 VSS VSS VCC VCC _0597_ sky130_fd_sc_hd__a21o_1
X_2553_ _0510_ _0526_ _0527_ VSS VSS VCC VCC _0528_ sky130_fd_sc_hd__o21ai_2
X_5341_ clknet_leaf_168_i_clk _0369_ VSS VSS VCC VCC u_muldiv.divisor\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_2484_ net647 net553 VSS VSS VCC VCC _0459_ sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_92_i_clk clknet_4_14__leaf_i_clk VSS VSS VCC VCC clknet_leaf_92_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5272_ clknet_4_10__leaf_i_clk _0300_ VSS VSS VCC VCC u_muldiv.quotient_msk\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_4223_ u_muldiv.divisor\[4\] _0444_ VSS VSS VCC VCC _1851_ sky130_fd_sc_hd__or2_2
X_4154_ net553 u_muldiv.i_on_wait net189 VSS VSS VCC VCC _0198_ sky130_fd_sc_hd__o21a_1
X_3105_ net445 net655 VSS VSS VCC VCC _1066_ sky130_fd_sc_hd__and2_1
X_4085_ net588 net587 VSS VSS VCC VCC _1794_ sky130_fd_sc_hd__or2_2
X_3036_ _0963_ _0969_ _0999_ _0965_ VSS VSS VCC VCC _1001_ sky130_fd_sc_hd__o211ai_4
Xclkbuf_leaf_30_i_clk clknet_4_4__leaf_i_clk VSS VSS VCC VCC clknet_leaf_30_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4987_ clknet_leaf_175_i_clk _0020_ VSS VSS VCC VCC u_bits.i_op1\[17\] sky130_fd_sc_hd__dfxtp_4
X_3938_ net233 net137 net396 VSS VSS VCC VCC _0101_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_45_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3869_ net506 net90 net719 VSS VSS VCC VCC _1684_ sky130_fd_sc_hd__a21o_1
Xfanout320 net321 VSS VSS VCC VCC net320 sky130_fd_sc_hd__buf_4
Xfanout331 _1722_ VSS VSS VCC VCC net331 sky130_fd_sc_hd__buf_6
Xfanout342 net343 VSS VSS VCC VCC net342 sky130_fd_sc_hd__buf_4
Xfanout353 _0783_ VSS VSS VCC VCC net353 sky130_fd_sc_hd__buf_2
Xfanout364 net365 VSS VSS VCC VCC net364 sky130_fd_sc_hd__clkbuf_8
Xfanout375 net376 VSS VSS VCC VCC net375 sky130_fd_sc_hd__buf_4
Xfanout386 net387 VSS VSS VCC VCC net386 sky130_fd_sc_hd__buf_4
Xfanout397 net398 VSS VSS VCC VCC net397 sky130_fd_sc_hd__buf_4
Xinput17 i_csr_data[1] VSS VSS VCC VCC net17 sky130_fd_sc_hd__buf_2
Xinput28 i_csr_data[2] VSS VSS VCC VCC net28 sky130_fd_sc_hd__clkbuf_4
Xinput39 i_flush VSS VSS VCC VCC net39 sky130_fd_sc_hd__buf_8
X_4910_ u_muldiv.divisor\[17\] net488 net341 u_muldiv.divisor\[18\] vssd1 vssd1 vccd1
+ vccd1 _0362_ sky130_fd_sc_hd__a22o_1
X_4841_ net660 _2368_ net369 net658 VSS VSS VCC VCC _2381_ sky130_fd_sc_hd__o211ai_1
X_4772_ _2316_ net371 net672 VSS VSS VCC VCC _2318_ sky130_fd_sc_hd__a21oi_1
X_3723_ net674 u_bits.i_op2\[21\] net412 _1599_ VSS VSS VCC VCC _1600_ sky130_fd_sc_hd__a31o_1
X_3654_ net607 _1280_ _0899_ _0856_ net409 VSS VSS VCC VCC _1536_ sky130_fd_sc_hd__a221o_1
X_2605_ _0534_ _0535_ _0542_ _0543_ VSS VSS VCC VCC _0580_ sky130_fd_sc_hd__o211ai_4
X_3585_ _1469_ _1470_ _1471_ VSS VSS VCC VCC _1472_ sky130_fd_sc_hd__o21ai_1
X_5324_ clknet_leaf_122_i_clk _0352_ VSS VSS VCC VCC u_muldiv.divisor\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2536_ net535 _0429_ VSS VSS VCC VCC _0511_ sky130_fd_sc_hd__nor2_1
X_5255_ clknet_leaf_94_i_clk _0283_ VSS VSS VCC VCC u_muldiv.quotient_msk\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2467_ net463 VSS VSS VCC VCC _0442_ sky130_fd_sc_hd__inv_2
X_4206_ op_cnt\[0\] op_cnt\[1\] op_cnt\[2\] VSS VSS VCC VCC _1838_ sky130_fd_sc_hd__and3_1
X_5186_ clknet_leaf_98_i_clk _0218_ VSS VSS VCC VCC u_muldiv.mul\[3\] sky130_fd_sc_hd__dfxtp_1
X_4137_ net580 _1831_ net570 VSS VSS VCC VCC _1835_ sky130_fd_sc_hd__o21bai_1
X_4068_ _1780_ net381 net590 VSS VSS VCC VCC _1781_ sky130_fd_sc_hd__a21oi_1
X_3019_ net661 u_bits.i_op2\[26\] _0984_ net348 VSS VSS VCC VCC _0985_ sky130_fd_sc_hd__o211a_1
X_3370_ _0781_ _1251_ _1240_ _1267_ VSS VSS VCC VCC _1268_ sky130_fd_sc_hd__o22ai_1
X_5040_ clknet_leaf_44_i_clk _0073_ VSS VSS VCC VCC u_bits.i_op2\[29\] sky130_fd_sc_hd__dfxtp_1
X_4824_ _1944_ _1946_ _1947_ VSS VSS VCC VCC _2365_ sky130_fd_sc_hd__nand3_1
X_4755_ _1720_ _2296_ _2302_ net317 VSS VSS VCC VCC _2303_ sky130_fd_sc_hd__o211ai_1
X_3706_ net613 _1044_ net607 VSS VSS VCC VCC _1584_ sky130_fd_sc_hd__o21a_1
X_4686_ _2222_ u_muldiv.dividend\[13\] net436 VSS VSS VCC VCC _2240_ sky130_fd_sc_hd__a21oi_1
X_3637_ u_bits.i_op2\[15\] net687 _1519_ net351 VSS VSS VCC VCC _1520_ sky130_fd_sc_hd__o211ai_1
X_3568_ _0976_ net606 _0766_ _1454_ VSS VSS VCC VCC _1456_ sky130_fd_sc_hd__a211o_2
X_5307_ clknet_4_2__leaf_i_clk _0335_ VSS VSS VCC VCC u_muldiv.dividend\[22\]
+ sky130_fd_sc_hd__dfxtp_2
X_2519_ net536 u_muldiv.add_prev\[19\] VSS VSS VCC VCC _0494_ sky130_fd_sc_hd__and2_1
X_3499_ _1391_ _1390_ _1388_ net443 VSS VSS VCC VCC _1392_ sky130_fd_sc_hd__a22o_2
X_5238_ clknet_leaf_126_i_clk _0266_ VSS VSS VCC VCC u_muldiv.o_div\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_5169_ clknet_leaf_70_i_clk _0201_ VSS VSS VCC VCC u_muldiv.add_prev\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_2870_ _0840_ net456 net651 _0767_ VSS VSS VCC VCC _0842_ sky130_fd_sc_hd__a31o_2
X_4540_ u_muldiv.quotient_msk\[28\] net477 net333 u_muldiv.quotient_msk\[29\] vssd1
+ vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__a22o_1
X_4471_ u_muldiv.o_div\[22\] _2077_ net319 VSS VSS VCC VCC _0273_ sky130_fd_sc_hd__mux2_1
X_3422_ net706 net704 net701 net700 net644 net633 VSS VSS VCC VCC _1318_ sky130_fd_sc_hd__mux4_1
X_3353_ u_wr_mux.i_reg_data2\[10\] _0764_ _1260_ VSS VSS VCC VCC net297 sky130_fd_sc_hd__a21o_4
X_3284_ net210 _1215_ VSS VSS VCC VCC _1216_ sky130_fd_sc_hd__nor2_1
X_5023_ clknet_leaf_49_i_clk _0056_ VSS VSS VCC VCC u_bits.i_op2\[12\] sky130_fd_sc_hd__dfxtp_2
X_4807_ net664 _2349_ VSS VSS VCC VCC _2350_ sky130_fd_sc_hd__nor2_1
X_2999_ _0965_ VSS VSS VCC VCC _0966_ sky130_fd_sc_hd__inv_2
X_4738_ _1917_ _2272_ _1909_ _1916_ VSS VSS VCC VCC _2287_ sky130_fd_sc_hd__o211a_1
X_4669_ _1895_ _1896_ _1892_ VSS VSS VCC VCC _2224_ sky130_fd_sc_hd__o21ai_1
X_3971_ u_wr_mux.i_reg_data2\[15\] net150 net397 VSS VSS VCC VCC _0133_ sky130_fd_sc_hd__mux2_1
X_2922_ net656 net654 net652 net651 net637 net625 VSS VSS VCC VCC _0892_ sky130_fd_sc_hd__mux4_2
X_2853_ net516 net523 _0823_ _0824_ VSS VSS VCC VCC _0826_ sky130_fd_sc_hd__a2bb2o_1
X_2784_ net560 net570 VSS VSS VCC VCC _0758_ sky130_fd_sc_hd__or2_4
X_4523_ u_muldiv.quotient_msk\[11\] net492 net339 u_muldiv.quotient_msk\[12\] vssd1
+ vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__a22o_1
X_4454_ net436 u_muldiv.quotient_msk\[19\] VSS VSS VCC VCC _2064_ sky130_fd_sc_hd__and2_1
X_3405_ _1300_ _1301_ net620 VSS VSS VCC VCC _1302_ sky130_fd_sc_hd__mux2_1
Xfanout705 u_bits.i_op1\[7\] VSS VSS VCC VCC net705 sky130_fd_sc_hd__clkbuf_8
X_4385_ _2006_ u_muldiv.o_div\[5\] net496 net385 VSS VSS VCC VCC _2009_ sky130_fd_sc_hd__a31o_1
Xfanout716 u_bits.i_op1\[2\] VSS VSS VCC VCC net716 sky130_fd_sc_hd__buf_4
Xfanout727 _1608_ VSS VSS VCC VCC net727 sky130_fd_sc_hd__buf_4
X_3336_ u_wr_mux.i_reg_data2\[12\] net305 net418 VSS VSS VCC VCC net282 sky130_fd_sc_hd__mux2_2
X_3267_ _0742_ _0731_ _0531_ VSS VSS VCC VCC _1205_ sky130_fd_sc_hd__o21ai_1
X_5006_ clknet_leaf_21_i_clk _0039_ VSS VSS VCC VCC net237 sky130_fd_sc_hd__dfxtp_4
X_3198_ _1153_ _1152_ net207 net355 net527 VSS VSS VCC VCC _1154_ sky130_fd_sc_hd__a221o_1
Xoutput308 net308 VSS VSS VCC VCC o_wdata[7] sky130_fd_sc_hd__buf_2
X_4170_ _1138_ _1139_ net400 VSS VSS VCC VCC _0214_ sky130_fd_sc_hd__and3_1
X_3121_ net632 net454 _0847_ _1080_ VSS VSS VCC VCC _1081_ sky130_fd_sc_hd__o31a_1
X_3052_ _1013_ net616 _1015_ VSS VSS VCC VCC _1016_ sky130_fd_sc_hd__a21oi_1
X_3954_ net182 net506 VSS VSS VCC VCC _1717_ sky130_fd_sc_hd__nand2b_1
X_2905_ _0874_ _0875_ VSS VSS VCC VCC _0876_ sky130_fd_sc_hd__nand2_1
X_3885_ net506 net94 net719 VSS VSS VCC VCC _1696_ sky130_fd_sc_hd__a21o_1
X_2836_ net679 net682 net684 net686 net637 net627 VSS VSS VCC VCC _0810_ sky130_fd_sc_hd__mux4_1
X_2767_ _0736_ _0685_ _0740_ VSS VSS VCC VCC _0742_ sky130_fd_sc_hd__a21o_2
X_4506_ _1990_ _1991_ _2102_ _2103_ _2104_ VSS VSS VCC VCC _2105_ sky130_fd_sc_hd__a221o_1
X_2698_ net445 u_bits.i_op2\[14\] VSS VSS VCC VCC _0673_ sky130_fd_sc_hd__nand2_1
X_4437_ _2042_ _0455_ VSS VSS VCC VCC _2050_ sky130_fd_sc_hd__nand2_4
Xfanout502 net503 VSS VSS VCC VCC net502 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout513 net514 VSS VSS VCC VCC net513 sky130_fd_sc_hd__clkbuf_2
Xfanout524 alu_ctrl\[2\] VSS VSS VCC VCC net524 sky130_fd_sc_hd__clkbuf_8
X_4368_ u_muldiv.quotient_msk\[1\] u_muldiv.o_div\[1\] net473 net438 vssd1 vssd1 vccd1
+ vccd1 _1996_ sky130_fd_sc_hd__o211a_1
Xfanout535 net536 VSS VSS VCC VCC net535 sky130_fd_sc_hd__buf_4
Xfanout546 net547 VSS VSS VCC VCC net546 sky130_fd_sc_hd__clkbuf_4
Xfanout557 net558 VSS VSS VCC VCC net557 sky130_fd_sc_hd__clkbuf_4
X_3319_ u_adder.i_cmp_inverse _1248_ VSS VSS VCC VCC _1249_ sky130_fd_sc_hd__nand2_1
Xfanout568 net569 VSS VSS VCC VCC net568 sky130_fd_sc_hd__buf_4
Xfanout579 u_bits.i_op2\[31\] VSS VSS VCC VCC net579 sky130_fd_sc_hd__buf_6
X_4299_ u_muldiv.dividend\[22\] u_muldiv.divisor\[22\] VSS VSS VCC VCC _1927_
+ sky130_fd_sc_hd__and2b_1
X_3670_ net589 net683 net349 _1550_ VSS VSS VCC VCC _1551_ sky130_fd_sc_hd__o211a_1
X_2621_ net539 _0425_ net431 _0594_ VSS VSS VCC VCC _0596_ sky130_fd_sc_hd__o211ai_4
X_5340_ clknet_leaf_167_i_clk _0368_ VSS VSS VCC VCC u_muldiv.divisor\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_2552_ _0498_ _0504_ _0505_ _0496_ VSS VSS VCC VCC _0527_ sky130_fd_sc_hd__a31oi_2
X_5271_ clknet_leaf_130_i_clk _0299_ VSS VSS VCC VCC u_muldiv.quotient_msk\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_2483_ net516 net524 VSS VSS VCC VCC _0458_ sky130_fd_sc_hd__or2_1
X_4222_ _0444_ u_muldiv.divisor\[4\] VSS VSS VCC VCC _1850_ sky130_fd_sc_hd__nand2_2
X_4153_ _1202_ _1203_ net401 VSS VSS VCC VCC _0197_ sky130_fd_sc_hd__and3_1
X_3104_ net533 u_muldiv.add_prev\[29\] VSS VSS VCC VCC _1065_ sky130_fd_sc_hd__and2_1
X_4084_ u_muldiv.divisor\[50\] net485 net336 u_muldiv.divisor\[51\] _1793_ vssd1 vssd1
+ vccd1 vccd1 _0170_ sky130_fd_sc_hd__a221o_1
X_3035_ _0969_ _0965_ _0963_ _0999_ VSS VSS VCC VCC _1000_ sky130_fd_sc_hd__a211o_2
X_4986_ clknet_leaf_92_i_clk _0019_ VSS VSS VCC VCC u_bits.i_op1\[16\] sky130_fd_sc_hd__dfxtp_4
X_3937_ net232 net136 net397 VSS VSS VCC VCC _0100_ sky130_fd_sc_hd__mux2_1
X_3868_ net506 _1682_ VSS VSS VCC VCC _1683_ sky130_fd_sc_hd__and2b_1
X_2819_ _0419_ net715 _0792_ VSS VSS VCC VCC _0793_ sky130_fd_sc_hd__a21oi_1
X_3799_ net600 net618 net545 VSS VSS VCC VCC _1631_ sky130_fd_sc_hd__mux2_1
Xfanout321 _1993_ VSS VSS VCC VCC net321 sky130_fd_sc_hd__buf_4
Xfanout332 net333 VSS VSS VCC VCC net332 sky130_fd_sc_hd__buf_4
Xfanout343 net344 VSS VSS VCC VCC net343 sky130_fd_sc_hd__buf_2
Xfanout354 net355 VSS VSS VCC VCC net354 sky130_fd_sc_hd__buf_4
Xfanout365 _0755_ VSS VSS VCC VCC net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 net377 VSS VSS VCC VCC net376 sky130_fd_sc_hd__buf_4
Xfanout387 net388 VSS VSS VCC VCC net387 sky130_fd_sc_hd__buf_6
Xfanout398 net399 VSS VSS VCC VCC net398 sky130_fd_sc_hd__buf_4
Xinput18 i_csr_data[20] VSS VSS VCC VCC net18 sky130_fd_sc_hd__clkbuf_4
Xinput29 i_csr_data[30] VSS VSS VCC VCC net29 sky130_fd_sc_hd__clkbuf_2
X_4840_ net670 net672 _2316_ _2379_ VSS VSS VCC VCC _2380_ sky130_fd_sc_hd__or4b_1
X_4771_ _2316_ net371 net672 VSS VSS VCC VCC _2317_ sky130_fd_sc_hd__and3_1
X_3722_ net674 u_bits.i_op2\[21\] net351 _1598_ VSS VSS VCC VCC _1599_ sky130_fd_sc_hd__o211a_1
X_3653_ net608 _1272_ net328 VSS VSS VCC VCC _1535_ sky130_fd_sc_hd__o21a_1
X_2604_ _0561_ _0554_ _0560_ _0568_ _0578_ VSS VSS VCC VCC _0579_ sky130_fd_sc_hd__o2111ai_4
X_3584_ u_bits.i_op2\[11\] net696 _0781_ net441 VSS VSS VCC VCC _1471_ sky130_fd_sc_hd__a211o_1
X_5323_ clknet_leaf_114_i_clk _0351_ VSS VSS VCC VCC u_muldiv.divisor\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_2535_ _0497_ _0498_ _0506_ _0507_ VSS VSS VCC VCC _0510_ sky130_fd_sc_hd__nand4_2
X_5254_ clknet_leaf_7_i_clk _0282_ VSS VSS VCC VCC u_muldiv.o_div\[31\] sky130_fd_sc_hd__dfxtp_1
X_2466_ u_muldiv.dividend\[3\] VSS VSS VCC VCC _0441_ sky130_fd_sc_hd__clkinv_2
X_4205_ op_cnt\[0\] op_cnt\[1\] op_cnt\[2\] VSS VSS VCC VCC _1837_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_112_i_clk clknet_4_14__leaf_i_clk VSS VSS VCC VCC clknet_leaf_112_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5185_ clknet_leaf_98_i_clk _0217_ VSS VSS VCC VCC u_muldiv.mul\[2\] sky130_fd_sc_hd__dfxtp_1
X_4136_ u_muldiv.divisor\[61\] net482 net337 u_muldiv.divisor\[62\] _1834_ vssd1 vssd1
+ vccd1 vccd1 _0181_ sky130_fd_sc_hd__a221o_1
X_4067_ u_bits.i_op2\[12\] _1774_ net591 _1764_ VSS VSS VCC VCC _1780_ sky130_fd_sc_hd__or4_2
X_3018_ net561 u_bits.i_op2\[26\] net661 VSS VSS VCC VCC _0984_ sky130_fd_sc_hd__nand3b_1
Xclkbuf_leaf_127_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_127_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4969_ _1248_ _2436_ _2437_ VSS VSS VCC VCC _0411_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_91_i_clk clknet_4_14__leaf_i_clk VSS VSS VCC VCC clknet_leaf_91_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_44_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_44_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_59_i_clk clknet_4_7__leaf_i_clk VSS VSS VCC VCC clknet_leaf_59_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4823_ _0449_ net323 _2364_ VSS VSS VCC VCC _0338_ sky130_fd_sc_hd__a21oi_1
X_4754_ _2298_ net434 _2297_ _2300_ _2301_ VSS VSS VCC VCC _2302_ sky130_fd_sc_hd__o32a_1
X_3705_ u_muldiv.mul\[52\] net361 net360 u_muldiv.mul\[20\] VSS VSS VCC VCC
+ _1583_ sky130_fd_sc_hd__a22o_1
X_4685_ u_muldiv.dividend\[13\] u_muldiv.dividend\[12\] u_muldiv.dividend\[11\] _2201_
+ VSS VSS VCC VCC _2239_ sky130_fd_sc_hd__or4_2
X_3636_ net564 net687 net591 VSS VSS VCC VCC _1519_ sky130_fd_sc_hd__nand3b_1
X_3567_ net607 net409 _0979_ VSS VSS VCC VCC _1455_ sky130_fd_sc_hd__or3_1
X_5306_ clknet_leaf_161_i_clk _0334_ VSS VSS VCC VCC u_muldiv.dividend\[21\]
+ sky130_fd_sc_hd__dfxtp_2
X_2518_ net516 net524 _0490_ _0491_ VSS VSS VCC VCC _0493_ sky130_fd_sc_hd__o211ai_2
X_3498_ net558 u_muldiv.mul\[5\] net415 net529 VSS VSS VCC VCC _1391_ sky130_fd_sc_hd__o31a_1
X_5237_ clknet_leaf_127_i_clk _0265_ VSS VSS VCC VCC u_muldiv.o_div\[14\]
+ sky130_fd_sc_hd__dfxtp_4
X_2449_ net733 VSS VSS VCC VCC _0424_ sky130_fd_sc_hd__inv_2
X_5168_ clknet_leaf_61_i_clk _0200_ VSS VSS VCC VCC u_muldiv.add_prev\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_4119_ net583 net382 _1817_ net582 VSS VSS VCC VCC _1821_ sky130_fd_sc_hd__a211o_1
X_5099_ clknet_leaf_172_i_clk _0132_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_4470_ _2075_ net488 _2074_ _2076_ VSS VSS VCC VCC _2077_ sky130_fd_sc_hd__a31o_1
X_3421_ net689 net687 net685 net683 net644 net632 VSS VSS VCC VCC _1317_ sky130_fd_sc_hd__mux4_2
X_3352_ net564 u_wr_mux.i_reg_data2\[26\] net417 net301 VSS VSS VCC VCC _1260_
+ sky130_fd_sc_hd__a22o_1
X_3283_ net208 _1214_ _1170_ _1165_ VSS VSS VCC VCC _1215_ sky130_fd_sc_hd__nand4b_1
X_5022_ clknet_leaf_15_i_clk _0055_ VSS VSS VCC VCC u_bits.i_op2\[11\] sky130_fd_sc_hd__dfxtp_4
X_4806_ net670 net672 net667 _2316_ net369 VSS VSS VCC VCC _2349_ sky130_fd_sc_hd__o41a_1
X_2998_ _0960_ _0961_ _0962_ VSS VSS VCC VCC _0965_ sky130_fd_sc_hd__nand3_4
X_4737_ _1909_ _1917_ _2273_ VSS VSS VCC VCC _2286_ sky130_fd_sc_hd__or3b_1
X_4668_ _2221_ _2222_ net437 VSS VSS VCC VCC _2223_ sky130_fd_sc_hd__a21o_1
X_3619_ net528 _1500_ _1502_ _1503_ VSS VSS VCC VCC _1504_ sky130_fd_sc_hd__a2bb2o_1
X_4599_ u_muldiv.dividend\[5\] _2147_ u_muldiv.dividend\[6\] VSS VSS VCC VCC
+ _2160_ sky130_fd_sc_hd__o21ai_1
X_3970_ u_wr_mux.i_reg_data2\[14\] net149 net386 VSS VSS VCC VCC _0132_ sky130_fd_sc_hd__mux2_1
X_2921_ net665 net662 net660 net658 net637 net625 VSS VSS VCC VCC _0891_ sky130_fd_sc_hd__mux4_2
X_2852_ _0823_ _0824_ net432 VSS VSS VCC VCC _0825_ sky130_fd_sc_hd__nand3_1
X_2783_ net562 net570 VSS VSS VCC VCC _0757_ sky130_fd_sc_hd__nor2_2
X_4522_ u_muldiv.quotient_msk\[10\] net492 net339 u_muldiv.quotient_msk\[11\] vssd1
+ vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__a22o_1
X_4453_ u_muldiv.o_div\[19\] _2060_ net470 net490 VSS VSS VCC VCC _2063_ sky130_fd_sc_hd__o2bb2a_1
X_3404_ net708 net706 net704 net701 net642 net628 VSS VSS VCC VCC _1301_ sky130_fd_sc_hd__mux4_1
X_4384_ u_muldiv.o_div\[4\] net331 net376 net320 _2008_ VSS VSS VCC VCC _0255_
+ sky130_fd_sc_hd__a32o_1
Xfanout706 u_bits.i_op1\[6\] VSS VSS VCC VCC net706 sky130_fd_sc_hd__buf_4
Xfanout717 net718 VSS VSS VCC VCC net717 sky130_fd_sc_hd__buf_6
Xfanout728 _1608_ VSS VSS VCC VCC net728 sky130_fd_sc_hd__clkbuf_4
X_3335_ u_wr_mux.i_reg_data2\[11\] net304 net416 VSS VSS VCC VCC net281 sky130_fd_sc_hd__mux2_8
X_3266_ _1204_ VSS VSS VCC VCC net188 sky130_fd_sc_hd__clkinv_4
X_5005_ clknet_leaf_31_i_clk _0038_ VSS VSS VCC VCC net236 sky130_fd_sc_hd__dfxtp_4
X_3197_ net411 _1146_ net522 VSS VSS VCC VCC _1153_ sky130_fd_sc_hd__a21oi_1
Xoutput309 net309 VSS VSS VCC VCC o_wdata[8] sky130_fd_sc_hd__buf_2
X_3120_ _0937_ net455 VSS VSS VCC VCC _1080_ sky130_fd_sc_hd__nand2_1
X_3051_ net346 _1014_ _0858_ _0905_ _0909_ VSS VSS VCC VCC _1015_ sky130_fd_sc_hd__o221ai_1
X_3953_ u_mux.i_add_override net5 net392 VSS VSS VCC VCC _0116_ sky130_fd_sc_hd__mux2_1
X_2904_ _0872_ _0873_ VSS VSS VCC VCC _0875_ sky130_fd_sc_hd__nand2_1
X_3884_ net506 _1694_ VSS VSS VCC VCC _1695_ sky130_fd_sc_hd__and2b_1
X_2835_ net458 net685 _0808_ VSS VSS VCC VCC _0809_ sky130_fd_sc_hd__a21oi_1
X_2766_ _0736_ _0685_ _0740_ VSS VSS VCC VCC _0741_ sky130_fd_sc_hd__a21oi_2
X_4505_ u_muldiv.quotient_msk\[30\] u_muldiv.o_div\[30\] net466 net433 vssd1 vssd1
+ vccd1 vccd1 _2104_ sky130_fd_sc_hd__o211a_1
X_2697_ net647 net552 net689 net535 net423 VSS VSS VCC VCC _0672_ sky130_fd_sc_hd__o2111ai_4
X_4436_ net322 _2047_ _2049_ _0455_ VSS VSS VCC VCC _0266_ sky130_fd_sc_hd__a2bb2oi_1
Xfanout503 net504 VSS VSS VCC VCC net503 sky130_fd_sc_hd__clkbuf_4
Xfanout514 net515 VSS VSS VCC VCC net514 sky130_fd_sc_hd__dlymetal6s2s_1
X_4367_ u_muldiv.o_div\[0\] u_muldiv.o_div\[1\] VSS VSS VCC VCC _1995_ sky130_fd_sc_hd__nand2_1
Xfanout525 alu_ctrl\[2\] VSS VSS VCC VCC net525 sky130_fd_sc_hd__buf_6
Xfanout536 net543 VSS VSS VCC VCC net536 sky130_fd_sc_hd__buf_4
Xfanout547 u_muldiv.i_is_div VSS VSS VCC VCC net547 sky130_fd_sc_hd__buf_4
X_3318_ _1246_ _1109_ _1135_ VSS VSS VCC VCC _1248_ sky130_fd_sc_hd__o21ai_2
Xfanout558 net559 VSS VSS VCC VCC net558 sky130_fd_sc_hd__clkbuf_4
Xfanout569 net216 VSS VSS VCC VCC net569 sky130_fd_sc_hd__buf_4
X_4298_ u_muldiv.divisor\[22\] u_muldiv.dividend\[22\] VSS VSS VCC VCC _1926_
+ sky130_fd_sc_hd__and2b_1
X_3249_ _0636_ _0637_ _0728_ VSS VSS VCC VCC _1191_ sky130_fd_sc_hd__a21boi_2
Xclkbuf_4_15__f_i_clk clknet_2_3_0_i_clk VSS VSS VCC VCC clknet_4_15__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2620_ net449 u_bits.i_op2\[5\] VSS VSS VCC VCC _0595_ sky130_fd_sc_hd__nand2_1
X_2551_ _0518_ _0525_ _0519_ VSS VSS VCC VCC _0526_ sky130_fd_sc_hd__a21boi_1
X_5270_ clknet_leaf_130_i_clk _0298_ VSS VSS VCC VCC u_muldiv.quotient_msk\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_2482_ net517 net524 VSS VSS VCC VCC _0457_ sky130_fd_sc_hd__nor2_8
X_4221_ _1847_ _1848_ VSS VSS VCC VCC _1849_ sky130_fd_sc_hd__nor2_2
X_4152_ _1194_ _1195_ net401 VSS VSS VCC VCC _0196_ sky130_fd_sc_hd__and3_1
X_3103_ net445 net581 _0464_ net655 net427 VSS VSS VCC VCC _1064_ sky130_fd_sc_hd__a221o_1
X_4083_ net587 _1791_ _1792_ VSS VSS VCC VCC _1793_ sky130_fd_sc_hd__a21oi_1
X_3034_ _0997_ _0998_ VSS VSS VCC VCC _0999_ sky130_fd_sc_hd__nand2_1
X_4985_ clknet_leaf_81_i_clk _0018_ VSS VSS VCC VCC u_bits.i_op1\[15\] sky130_fd_sc_hd__dfxtp_1
X_3936_ net231 net135 net399 VSS VSS VCC VCC _0099_ sky130_fd_sc_hd__mux2_1
X_3867_ u_bits.i_op2\[22\] u_bits.i_op2\[20\] net547 VSS VSS VCC VCC _1682_
+ sky130_fd_sc_hd__mux2_1
X_2818_ net645 net717 VSS VSS VCC VCC _0792_ sky130_fd_sc_hd__and2_1
X_3798_ net618 net727 _1630_ _1629_ VSS VSS VCC VCC _0047_ sky130_fd_sc_hd__o22a_1
X_2749_ _0718_ _0719_ _0722_ _0723_ VSS VSS VCC VCC _0724_ sky130_fd_sc_hd__o2bb2ai_4
X_4419_ _2019_ _2034_ _0452_ _0453_ _0454_ VSS VSS VCC VCC _2036_ sky130_fd_sc_hd__a41o_1
Xfanout322 net323 VSS VSS VCC VCC net322 sky130_fd_sc_hd__buf_6
Xfanout333 net334 VSS VSS VCC VCC net333 sky130_fd_sc_hd__buf_6
Xfanout344 _1719_ VSS VSS VCC VCC net344 sky130_fd_sc_hd__buf_12
Xfanout355 _0763_ VSS VSS VCC VCC net355 sky130_fd_sc_hd__buf_6
Xfanout366 net367 VSS VSS VCC VCC net366 sky130_fd_sc_hd__buf_4
Xfanout377 _1991_ VSS VSS VCC VCC net377 sky130_fd_sc_hd__buf_8
Xfanout388 _1610_ VSS VSS VCC VCC net388 sky130_fd_sc_hd__buf_6
Xfanout399 _1610_ VSS VSS VCC VCC net399 sky130_fd_sc_hd__buf_2
Xinput19 i_csr_data[21] VSS VSS VCC VCC net19 sky130_fd_sc_hd__clkbuf_1
X_4770_ net679 net677 net675 _2290_ VSS VSS VCC VCC _2316_ sky130_fd_sc_hd__or4_4
X_3721_ net569 _0431_ net674 VSS VSS VCC VCC _1598_ sky130_fd_sc_hd__or3b_1
X_3652_ u_muldiv.mul\[48\] net361 net360 u_muldiv.mul\[16\] VSS VSS VCC VCC
+ _1534_ sky130_fd_sc_hd__a22oi_1
X_2603_ _0569_ _0577_ VSS VSS VCC VCC _0578_ sky130_fd_sc_hd__nand2_2
X_3583_ net572 net421 _1011_ net345 _1466_ VSS VSS VCC VCC _1470_ sky130_fd_sc_hd__a221o_1
X_2534_ _0508_ VSS VSS VCC VCC _0509_ sky130_fd_sc_hd__clkinv_2
X_5322_ clknet_leaf_115_i_clk _0350_ VSS VSS VCC VCC u_muldiv.divisor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2465_ u_muldiv.dividend\[0\] VSS VSS VCC VCC _0440_ sky130_fd_sc_hd__inv_2
X_5253_ clknet_leaf_7_i_clk _0281_ VSS VSS VCC VCC u_muldiv.o_div\[30\] sky130_fd_sc_hd__dfxtp_2
X_4204_ op_cnt\[0\] op_cnt\[1\] _1836_ VSS VSS VCC VCC _0247_ sky130_fd_sc_hd__o21a_1
X_5184_ clknet_leaf_104_i_clk _0216_ VSS VSS VCC VCC u_muldiv.mul\[1\] sky130_fd_sc_hd__dfxtp_1
X_4135_ _1832_ _1833_ VSS VSS VCC VCC _1834_ sky130_fd_sc_hd__nor2_1
X_4066_ u_bits.i_op2\[12\] _1774_ net591 _1764_ VSS VSS VCC VCC _1779_ sky130_fd_sc_hd__nor4_1
X_3017_ _0982_ net346 net450 _0980_ _0981_ VSS VSS VCC VCC _0983_ sky130_fd_sc_hd__o221a_1
X_4968_ _1248_ _2436_ net400 VSS VSS VCC VCC _2437_ sky130_fd_sc_hd__a21oi_1
X_3919_ u_pc_sel.i_pc_next\[10\] net109 net394 VSS VSS VCC VCC _0085_ sky130_fd_sc_hd__mux2_1
X_4899_ u_muldiv.divisor\[6\] net493 net339 u_muldiv.divisor\[7\] vssd1 vssd1 vccd1
+ vccd1 _0351_ sky130_fd_sc_hd__a22o_1
X_4822_ _2357_ _2361_ _2363_ net315 VSS VSS VCC VCC _2364_ sky130_fd_sc_hd__o211a_1
X_4753_ net677 _2299_ net481 net467 VSS VSS VCC VCC _2301_ sky130_fd_sc_hd__a211o_1
X_3704_ u_muldiv.dividend\[20\] net420 net368 u_muldiv.o_div\[20\] vssd1 vssd1 vccd1
+ vccd1 _1582_ sky130_fd_sc_hd__a22o_1
X_4684_ _2233_ _2232_ _2237_ VSS VSS VCC VCC _2238_ sky130_fd_sc_hd__a21oi_1
X_3635_ net574 u_pc_sel.i_pc_next\[14\] _1517_ _1518_ VSS VSS VCC VCC net250
+ sky130_fd_sc_hd__a22o_4
X_3566_ net606 _1453_ VSS VSS VCC VCC _1454_ sky130_fd_sc_hd__nor2_1
X_5305_ clknet_leaf_160_i_clk _0333_ VSS VSS VCC VCC u_muldiv.dividend\[20\]
+ sky130_fd_sc_hd__dfxtp_2
X_2517_ _0490_ _0491_ net516 net523 VSS VSS VCC VCC _0492_ sky130_fd_sc_hd__a211o_1
X_3497_ net441 u_muldiv.mul\[37\] net414 _1389_ VSS VSS VCC VCC _1390_ sky130_fd_sc_hd__a31o_1
X_2448_ net541 VSS VSS VCC VCC _0423_ sky130_fd_sc_hd__inv_4
X_5236_ clknet_leaf_127_i_clk _0264_ VSS VSS VCC VCC u_muldiv.o_div\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_5167_ clknet_leaf_74_i_clk _0199_ VSS VSS VCC VCC u_muldiv.add_prev\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_4118_ net583 _1816_ net382 net582 VSS VSS VCC VCC _1820_ sky130_fd_sc_hd__o211ai_1
X_5098_ clknet_leaf_175_i_clk _0131_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[13\]
+ sky130_fd_sc_hd__dfxtp_4
X_4049_ _1764_ net381 net593 net330 VSS VSS VCC VCC _1766_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_173_i_clk clknet_4_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_173_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_4_3__f_i_clk clknet_2_0_0_i_clk VSS VSS VCC VCC clknet_4_3__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_111_i_clk clknet_4_9__leaf_i_clk VSS VSS VCC VCC clknet_leaf_111_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3420_ net697 net696 net694 net692 net645 net633 VSS VSS VCC VCC _1316_ sky130_fd_sc_hd__mux4_2
Xclkbuf_leaf_126_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_126_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3351_ u_wr_mux.i_reg_data2\[9\] _0764_ _1259_ VSS VSS VCC VCC net296 sky130_fd_sc_hd__a21o_1
X_3282_ _0576_ _1211_ net194 VSS VSS VCC VCC _1214_ sky130_fd_sc_hd__a21oi_4
X_5021_ clknet_leaf_14_i_clk _0054_ VSS VSS VCC VCC u_bits.i_op2\[10\] sky130_fd_sc_hd__dfxtp_4
X_4805_ _1946_ _1944_ net466 VSS VSS VCC VCC _2348_ sky130_fd_sc_hd__o21ai_1
X_2997_ _0960_ _0961_ _0962_ VSS VSS VCC VCC _0964_ sky130_fd_sc_hd__a21o_1
X_4736_ _2283_ _2284_ net437 VSS VSS VCC VCC _2285_ sky130_fd_sc_hd__a21oi_1
X_4667_ u_muldiv.dividend\[11\] _2194_ _0446_ _0445_ VSS VSS VCC VCC _2222_
+ sky130_fd_sc_hd__nand4b_4
X_3618_ net557 u_muldiv.mul\[13\] net413 net528 VSS VSS VCC VCC _1503_ sky130_fd_sc_hd__o31a_1
X_4598_ u_muldiv.dividend\[5\] net325 net376 _2159_ VSS VSS VCC VCC _0318_
+ sky130_fd_sc_hd__a31o_1
X_3549_ _0934_ net604 VSS VSS VCC VCC _1438_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_leaf_90_i_clk clknet_4_15__leaf_i_clk VSS VSS VCC VCC clknet_leaf_90_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_5219_ clknet_leaf_45_i_clk _0248_ VSS VSS VCC VCC op_cnt\[2\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_43_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_43_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_58_i_clk clknet_4_7__leaf_i_clk VSS VSS VCC VCC clknet_leaf_58_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2920_ net650 u_bits.i_sra net451 VSS VSS VCC VCC _0890_ sky130_fd_sc_hd__a21o_1
X_2851_ net446 u_bits.i_op2\[23\] VSS VSS VCC VCC _0824_ sky130_fd_sc_hd__nand2_1
X_2782_ u_muldiv.dividend\[22\] net419 net365 u_muldiv.o_div\[22\] net442 vssd1 vssd1
+ vccd1 vccd1 _0756_ sky130_fd_sc_hd__a221o_1
X_4521_ u_muldiv.quotient_msk\[9\] net492 net339 u_muldiv.quotient_msk\[10\] vssd1
+ vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__a22o_1
X_4452_ net322 _2062_ _1998_ u_muldiv.o_div\[18\] VSS VSS VCC VCC _0269_ sky130_fd_sc_hd__a2bb2o_1
X_3403_ net717 net715 net713 net710 net642 net628 VSS VSS VCC VCC _1300_ sky130_fd_sc_hd__mux4_1
X_4383_ _2006_ _2007_ net496 net342 u_muldiv.quotient_msk\[4\] VSS VSS VCC VCC
+ _2008_ sky130_fd_sc_hd__a32o_1
Xfanout707 u_bits.i_op1\[6\] VSS VSS VCC VCC net707 sky130_fd_sc_hd__buf_4
X_3334_ u_wr_mux.i_reg_data2\[10\] net301 net417 VSS VSS VCC VCC net280 sky130_fd_sc_hd__mux2_4
Xfanout718 u_bits.i_op1\[1\] VSS VSS VCC VCC net718 sky130_fd_sc_hd__buf_4
Xfanout729 net730 VSS VSS VCC VCC net729 sky130_fd_sc_hd__buf_8
X_3265_ _1202_ _1203_ VSS VSS VCC VCC _1204_ sky130_fd_sc_hd__nand2_4
X_5004_ clknet_leaf_58_i_clk _0037_ VSS VSS VCC VCC net235 sky130_fd_sc_hd__dfxtp_4
X_3196_ _0909_ _1145_ _1149_ _1151_ VSS VSS VCC VCC _1152_ sky130_fd_sc_hd__a211o_1
X_4719_ _0413_ _2268_ _2269_ net488 VSS VSS VCC VCC _2270_ sky130_fd_sc_hd__a31o_1
X_3050_ net659 net661 net663 net666 net639 net636 VSS VSS VCC VCC _1014_ sky130_fd_sc_hd__mux4_1
X_3952_ u_bits.i_sra net4 net387 VSS VSS VCC VCC _0115_ sky130_fd_sc_hd__mux2_1
X_2903_ _0873_ _0872_ VSS VSS VCC VCC _0874_ sky130_fd_sc_hd__or2_1
X_3883_ net583 net585 net545 VSS VSS VCC VCC _1694_ sky130_fd_sc_hd__mux2_1
X_2834_ net643 net686 VSS VSS VCC VCC _0808_ sky130_fd_sc_hd__and2_1
X_2765_ _0684_ _0738_ _0739_ _0669_ VSS VSS VCC VCC _0740_ sky130_fd_sc_hd__o211ai_2
X_4504_ u_muldiv.o_div\[28\] u_muldiv.o_div\[29\] u_muldiv.o_div\[30\] _2094_ net477
+ VSS VSS VCC VCC _2103_ sky130_fd_sc_hd__o41a_1
X_2696_ _0669_ _0670_ VSS VSS VCC VCC _0671_ sky130_fd_sc_hd__nand2_2
X_4435_ net324 net376 _2043_ _2048_ VSS VSS VCC VCC _2049_ sky130_fd_sc_hd__a22o_1
Xfanout504 net240 VSS VSS VCC VCC net504 sky130_fd_sc_hd__clkbuf_4
Xfanout515 net240 VSS VSS VCC VCC net515 sky130_fd_sc_hd__clkbuf_2
X_4366_ u_muldiv.o_div\[0\] u_muldiv.o_div\[1\] VSS VSS VCC VCC _1994_ sky130_fd_sc_hd__or2_1
Xfanout526 alu_ctrl\[2\] VSS VSS VCC VCC net526 sky130_fd_sc_hd__clkbuf_4
Xfanout537 net539 VSS VSS VCC VCC net537 sky130_fd_sc_hd__clkbuf_4
Xfanout548 net550 VSS VSS VCC VCC net548 sky130_fd_sc_hd__buf_4
X_3317_ _1108_ _1101_ _1106_ _1136_ VSS VSS VCC VCC _1247_ sky130_fd_sc_hd__o211a_1
Xfanout559 net217 VSS VSS VCC VCC net559 sky130_fd_sc_hd__buf_6
X_4297_ _1908_ _1920_ _1924_ VSS VSS VCC VCC _1925_ sky130_fd_sc_hd__a21oi_4
X_3248_ _1190_ VSS VSS VCC VCC net184 sky130_fd_sc_hd__clkinv_4
X_3179_ _1133_ _1134_ _1128_ VSS VSS VCC VCC _1136_ sky130_fd_sc_hd__a21bo_1
X_2550_ _0522_ _0523_ _0524_ VSS VSS VCC VCC _0525_ sky130_fd_sc_hd__a21boi_4
X_2481_ u_muldiv.o_div\[20\] VSS VSS VCC VCC _0456_ sky130_fd_sc_hd__inv_2
X_4220_ u_muldiv.dividend\[5\] u_muldiv.divisor\[5\] VSS VSS VCC VCC _1848_
+ sky130_fd_sc_hd__and2b_1
X_4151_ _1193_ _1197_ net401 VSS VSS VCC VCC _0195_ sky130_fd_sc_hd__and3_1
X_3102_ net516 net524 _1062_ VSS VSS VCC VCC _1063_ sky130_fd_sc_hd__o21ai_1
X_4082_ net587 _1791_ net384 VSS VSS VCC VCC _1792_ sky130_fd_sc_hd__o21ai_1
X_3033_ _0993_ _0994_ _0995_ VSS VSS VCC VCC _0998_ sky130_fd_sc_hd__a21o_1
X_4984_ clknet_leaf_143_i_clk _0017_ VSS VSS VCC VCC u_bits.i_op1\[14\] sky130_fd_sc_hd__dfxtp_1
X_3935_ net230 net134 net386 VSS VSS VCC VCC _0098_ sky130_fd_sc_hd__mux2_1
X_3866_ u_bits.i_op2\[20\] net723 _1681_ _1680_ VSS VSS VCC VCC _0064_ sky130_fd_sc_hd__o22a_1
X_2817_ net458 net460 VSS VSS VCC VCC _0791_ sky130_fd_sc_hd__nand2_1
X_3797_ net511 net102 net721 VSS VSS VCC VCC _1630_ sky130_fd_sc_hd__a21o_1
X_2748_ u_muldiv.add_prev\[9\] net448 VSS VSS VCC VCC _0723_ sky130_fd_sc_hd__nor2_1
X_2679_ net519 net525 net592 net448 VSS VSS VCC VCC _0654_ sky130_fd_sc_hd__a2bb2o_1
X_4418_ _2027_ _2034_ _0454_ VSS VSS VCC VCC _2035_ sky130_fd_sc_hd__nand3_4
Xfanout323 _1992_ VSS VSS VCC VCC net323 sky130_fd_sc_hd__buf_12
Xfanout334 net344 VSS VSS VCC VCC net334 sky130_fd_sc_hd__buf_6
X_4349_ u_muldiv.divisor\[51\] u_muldiv.divisor\[50\] u_muldiv.divisor\[49\] u_muldiv.divisor\[48\]
+ VSS VSS VCC VCC _1977_ sky130_fd_sc_hd__or4_4
Xfanout345 _0909_ VSS VSS VCC VCC net345 sky130_fd_sc_hd__buf_4
Xfanout356 _0762_ VSS VSS VCC VCC net356 sky130_fd_sc_hd__buf_6
Xfanout367 net368 VSS VSS VCC VCC net367 sky130_fd_sc_hd__clkbuf_4
Xfanout378 net382 VSS VSS VCC VCC net378 sky130_fd_sc_hd__clkbuf_4
Xfanout389 net390 VSS VSS VCC VCC net389 sky130_fd_sc_hd__buf_4
X_3720_ net605 _1380_ net327 VSS VSS VCC VCC _1597_ sky130_fd_sc_hd__o21a_1
X_3651_ u_muldiv.dividend\[16\] net420 net368 u_muldiv.o_div\[16\] vssd1 vssd1 vccd1
+ vccd1 _1533_ sky130_fd_sc_hd__a22oi_1
X_2602_ net431 _0573_ _0576_ VSS VSS VCC VCC _0577_ sky130_fd_sc_hd__o21a_2
X_3582_ net608 _1468_ _0765_ _1467_ VSS VSS VCC VCC _1469_ sky130_fd_sc_hd__o211a_1
X_5321_ clknet_leaf_93_i_clk _0349_ VSS VSS VCC VCC u_muldiv.divisor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2533_ _0506_ _0507_ VSS VSS VCC VCC _0508_ sky130_fd_sc_hd__nand2_1
X_5252_ clknet_leaf_7_i_clk _0280_ VSS VSS VCC VCC u_muldiv.o_div\[29\] sky130_fd_sc_hd__dfxtp_2
X_2464_ net693 VSS VSS VCC VCC _0439_ sky130_fd_sc_hd__inv_2
X_4203_ op_cnt\[0\] op_cnt\[1\] net509 VSS VSS VCC VCC _1836_ sky130_fd_sc_hd__a21oi_1
X_5183_ clknet_leaf_104_i_clk _0215_ VSS VSS VCC VCC u_muldiv.mul\[0\] sky130_fd_sc_hd__dfxtp_1
X_4134_ _1831_ net378 net580 net330 VSS VSS VCC VCC _1833_ sky130_fd_sc_hd__a31o_1
X_4065_ u_muldiv.divisor\[46\] net485 net336 u_muldiv.divisor\[47\] _1778_ vssd1 vssd1
+ vccd1 vccd1 _0166_ sky130_fd_sc_hd__a221o_1
X_3016_ net660 net663 net664 net667 net638 net627 VSS VSS VCC VCC _0982_ sky130_fd_sc_hd__mux4_1
X_4967_ net517 _0781_ VSS VSS VCC VCC _2436_ sky130_fd_sc_hd__nor2_1
X_3918_ u_pc_sel.i_pc_next\[9\] net123 net386 VSS VSS VCC VCC _0084_ sky130_fd_sc_hd__mux2_1
X_4898_ u_muldiv.divisor\[5\] net496 net342 u_muldiv.divisor\[6\] vssd1 vssd1 vccd1
+ vccd1 _0350_ sky130_fd_sc_hd__a22o_1
X_3849_ net508 net84 net722 VSS VSS VCC VCC _1669_ sky130_fd_sc_hd__a21o_1
X_4821_ u_muldiv.dividend\[25\] _2345_ _2362_ VSS VSS VCC VCC _2363_ sky130_fd_sc_hd__o21ai_1
X_4752_ net677 _2299_ VSS VSS VCC VCC _2300_ sky130_fd_sc_hd__nor2_1
X_3703_ net729 net16 _1581_ VSS VSS VCC VCC net255 sky130_fd_sc_hd__o21a_4
X_4683_ net489 _2235_ _2236_ _1720_ VSS VSS VCC VCC _2237_ sky130_fd_sc_hd__o31a_1
X_3634_ net11 net730 net574 VSS VSS VCC VCC _1518_ sky130_fd_sc_hd__o21ba_1
X_3565_ _0770_ _1317_ _1319_ _1316_ net451 net456 VSS VSS VCC VCC _1453_ sky130_fd_sc_hd__mux4_1
X_5304_ clknet_leaf_148_i_clk _0332_ VSS VSS VCC VCC u_muldiv.dividend\[19\]
+ sky130_fd_sc_hd__dfxtp_4
X_2516_ net445 net587 VSS VSS VCC VCC _0491_ sky130_fd_sc_hd__nand2_1
X_3496_ u_muldiv.dividend\[5\] net420 net366 u_muldiv.o_div\[5\] net358 vssd1 vssd1
+ vccd1 vccd1 _1389_ sky130_fd_sc_hd__a221o_1
X_5235_ clknet_leaf_118_i_clk _0263_ VSS VSS VCC VCC u_muldiv.o_div\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_2447_ net521 VSS VSS VCC VCC _0422_ sky130_fd_sc_hd__inv_6
X_5166_ clknet_4_13__leaf_i_clk _0198_ VSS VSS VCC VCC u_muldiv.add_prev\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_4117_ u_muldiv.divisor\[57\] net483 net337 u_muldiv.divisor\[58\] _1819_ vssd1 vssd1
+ vccd1 vccd1 _0177_ sky130_fd_sc_hd__a221o_1
X_5097_ clknet_leaf_46_i_clk _0130_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[12\]
+ sky130_fd_sc_hd__dfxtp_4
X_4048_ _1764_ net381 net593 VSS VSS VCC VCC _1765_ sky130_fd_sc_hd__a21oi_1
Xoutput290 net290 VSS VSS VCC VCC o_wdata[1] sky130_fd_sc_hd__buf_2
X_3350_ net563 u_wr_mux.i_reg_data2\[25\] net416 net290 VSS VSS VCC VCC _1259_
+ sky130_fd_sc_hd__a22o_1
X_3281_ net194 VSS VSS VCC VCC _1213_ sky130_fd_sc_hd__clkinv_4
X_5020_ clknet_4_7__leaf_i_clk _0053_ VSS VSS VCC VCC u_bits.i_op2\[9\] sky130_fd_sc_hd__dfxtp_4
X_4804_ _1944_ _1946_ VSS VSS VCC VCC _2347_ sky130_fd_sc_hd__and2_1
X_2996_ _0960_ _0961_ _0962_ VSS VSS VCC VCC _0963_ sky130_fd_sc_hd__a21oi_2
X_4735_ u_muldiv.dividend\[18\] net462 u_muldiv.dividend\[16\] _2258_ vssd1 vssd1
+ vccd1 vccd1 _2284_ sky130_fd_sc_hd__or4_2
X_4666_ u_muldiv.dividend\[11\] _2201_ u_muldiv.dividend\[12\] VSS VSS VCC VCC
+ _2221_ sky130_fd_sc_hd__o21ai_1
X_3617_ _0434_ u_muldiv.mul\[45\] net413 _1501_ VSS VSS VCC VCC _1502_ sky130_fd_sc_hd__a31o_1
X_4597_ net325 net376 _2152_ _2158_ VSS VSS VCC VCC _2159_ sky130_fd_sc_hd__a211oi_1
X_3548_ net578 u_pc_sel.i_pc_next\[8\] _1436_ _1437_ VSS VSS VCC VCC net275
+ sky130_fd_sc_hd__a22o_2
X_3479_ _1372_ _1371_ net209 net354 VSS VSS VCC VCC _1373_ sky130_fd_sc_hd__a2bb2o_1
X_5218_ clknet_leaf_45_i_clk _0247_ VSS VSS VCC VCC op_cnt\[1\] sky130_fd_sc_hd__dfxtp_1
X_5149_ clknet_leaf_13_i_clk _0181_ VSS VSS VCC VCC u_muldiv.divisor\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_2850_ net641 net552 net669 net535 net424 VSS VSS VCC VCC _0823_ sky130_fd_sc_hd__o2111ai_1
X_2781_ net566 net441 VSS VSS VCC VCC _0755_ sky130_fd_sc_hd__nor2_4
X_4520_ u_muldiv.quotient_msk\[8\] net493 net339 u_muldiv.quotient_msk\[9\] vssd1
+ vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__a22o_1
X_4451_ u_muldiv.quotient_msk\[18\] net338 _2061_ _2060_ VSS VSS VCC VCC _2062_
+ sky130_fd_sc_hd__a22oi_1
X_3402_ _1297_ _1298_ net455 VSS VSS VCC VCC _1299_ sky130_fd_sc_hd__mux2_1
X_4382_ _2005_ u_muldiv.o_div\[4\] VSS VSS VCC VCC _2007_ sky130_fd_sc_hd__nand2_1
X_3333_ u_wr_mux.i_reg_data2\[9\] net290 net416 VSS VSS VCC VCC net310 sky130_fd_sc_hd__mux2_2
Xfanout708 u_bits.i_op1\[5\] VSS VSS VCC VCC net708 sky130_fd_sc_hd__buf_6
Xfanout719 net720 VSS VSS VCC VCC net719 sky130_fd_sc_hd__clkbuf_4
X_3264_ _0738_ _1199_ _0683_ VSS VSS VCC VCC _1203_ sky130_fd_sc_hd__a21o_1
X_5003_ clknet_leaf_30_i_clk _0036_ VSS VSS VCC VCC net241 sky130_fd_sc_hd__dfxtp_2
X_3195_ _0901_ _1150_ VSS VSS VCC VCC _1151_ sky130_fd_sc_hd__nor2_1
X_2979_ net673 net677 net675 net679 net627 net637 VSS VSS VCC VCC _0947_ sky130_fd_sc_hd__mux4_2
Xclkbuf_leaf_172_i_clk clknet_4_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_172_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4718_ _2266_ _2114_ net684 VSS VSS VCC VCC _2269_ sky130_fd_sc_hd__or3b_1
X_4649_ net701 net699 _2184_ VSS VSS VCC VCC _2206_ sky130_fd_sc_hd__nor3_2
Xclkbuf_leaf_110_i_clk clknet_4_11__leaf_i_clk VSS VSS VCC VCC clknet_leaf_110_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_125_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_125_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3951_ net526 net3 net399 VSS VSS VCC VCC _0114_ sky130_fd_sc_hd__mux2_1
X_2902_ net666 u_muldiv.add_prev\[24\] net534 VSS VSS VCC VCC _0873_ sky130_fd_sc_hd__mux2_1
X_3882_ net585 net724 _1693_ _1692_ VSS VSS VCC VCC _0068_ sky130_fd_sc_hd__o22a_1
X_2833_ net608 net616 VSS VSS VCC VCC _0807_ sky130_fd_sc_hd__or2_4
X_2764_ _0679_ _0670_ VSS VSS VCC VCC _0739_ sky130_fd_sc_hd__nand2_1
X_4503_ u_muldiv.o_div\[29\] _2095_ u_muldiv.o_div\[30\] VSS VSS VCC VCC _2102_
+ sky130_fd_sc_hd__o21ai_1
X_2695_ _0668_ _0666_ _0665_ VSS VSS VCC VCC _0670_ sky130_fd_sc_hd__nand3b_2
X_4434_ net436 u_muldiv.quotient_msk\[15\] VSS VSS VCC VCC _2048_ sky130_fd_sc_hd__nand2_1
X_4365_ net326 net377 VSS VSS VCC VCC _1993_ sky130_fd_sc_hd__nand2_8
Xfanout505 net506 VSS VSS VCC VCC net505 sky130_fd_sc_hd__buf_2
Xfanout516 net517 VSS VSS VCC VCC net516 sky130_fd_sc_hd__clkbuf_8
Xfanout527 net544 VSS VSS VCC VCC net527 sky130_fd_sc_hd__buf_8
Xfanout538 net539 VSS VSS VCC VCC net538 sky130_fd_sc_hd__buf_2
X_3316_ _1106_ _1136_ VSS VSS VCC VCC _1246_ sky130_fd_sc_hd__nand2_1
Xfanout549 net550 VSS VSS VCC VCC net549 sky130_fd_sc_hd__buf_4
X_4296_ _1923_ u_muldiv.divisor\[18\] _1910_ _1922_ VSS VSS VCC VCC _1924_
+ sky130_fd_sc_hd__o211ai_2
X_3247_ _1185_ _1189_ VSS VSS VCC VCC _1190_ sky130_fd_sc_hd__nand2_2
X_3178_ _1128_ _1133_ _1134_ VSS VSS VCC VCC _1135_ sky130_fd_sc_hd__nand3b_1
Xclkbuf_leaf_42_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_42_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2480_ u_muldiv.o_div\[15\] VSS VSS VCC VCC _0455_ sky130_fd_sc_hd__inv_2
X_4150_ _1186_ _1187_ net401 VSS VSS VCC VCC _0194_ sky130_fd_sc_hd__and3_1
X_3101_ net445 net581 _0464_ net655 VSS VSS VCC VCC _1062_ sky130_fd_sc_hd__a22o_1
X_4081_ net590 net589 u_bits.i_op2\[18\] _1780_ net380 VSS VSS VCC VCC _1791_
+ sky130_fd_sc_hd__o41a_1
X_3032_ _0993_ _0994_ _0995_ VSS VSS VCC VCC _0997_ sky130_fd_sc_hd__nand3_1
X_4983_ clknet_leaf_117_i_clk _0016_ VSS VSS VCC VCC u_bits.i_op1\[13\] sky130_fd_sc_hd__dfxtp_1
X_3934_ net229 net133 net393 VSS VSS VCC VCC _0097_ sky130_fd_sc_hd__mux2_1
X_3865_ net502 net89 net720 VSS VSS VCC VCC _1681_ sky130_fd_sc_hd__a21o_1
X_2816_ net649 _0435_ _0789_ VSS VSS VCC VCC _0790_ sky130_fd_sc_hd__o21a_1
X_3796_ net511 _1628_ VSS VSS VCC VCC _1629_ sky130_fd_sc_hd__and2b_1
X_2747_ net541 net700 VSS VSS VCC VCC _0722_ sky130_fd_sc_hd__nor2_1
X_2678_ net448 net592 VSS VSS VCC VCC _0653_ sky130_fd_sc_hd__nand2_1
X_4417_ u_muldiv.o_div\[10\] u_muldiv.o_div\[11\] VSS VSS VCC VCC _2034_ sky130_fd_sc_hd__nor2_1
X_4348_ u_muldiv.divisor\[61\] u_muldiv.divisor\[60\] u_muldiv.divisor\[62\] net482
+ VSS VSS VCC VCC _1976_ sky130_fd_sc_hd__or4_2
Xfanout324 net326 VSS VSS VCC VCC net324 sky130_fd_sc_hd__buf_4
Xfanout335 net337 VSS VSS VCC VCC net335 sky130_fd_sc_hd__clkbuf_4
Xfanout346 _0908_ VSS VSS VCC VCC net346 sky130_fd_sc_hd__buf_6
Xfanout357 _0760_ VSS VSS VCC VCC net357 sky130_fd_sc_hd__buf_4
Xfanout368 _0755_ VSS VSS VCC VCC net368 sky130_fd_sc_hd__buf_6
Xfanout379 net382 VSS VSS VCC VCC net379 sky130_fd_sc_hd__clkbuf_4
X_4279_ _0414_ _1904_ u_muldiv.dividend\[14\] _1903_ VSS VSS VCC VCC _1907_
+ sky130_fd_sc_hd__a31o_1
X_3650_ net576 u_pc_sel.i_pc_next\[15\] _1531_ _1532_ VSS VSS VCC VCC net251
+ sky130_fd_sc_hd__a22o_2
X_2601_ _0570_ _0572_ _0574_ _0575_ VSS VSS VCC VCC _0576_ sky130_fd_sc_hd__o2bb2ai_4
X_3581_ _0837_ _1337_ _1339_ _1340_ net457 net452 VSS VSS VCC VCC _1468_ sky130_fd_sc_hd__mux4_1
X_5320_ clknet_leaf_92_i_clk _0348_ VSS VSS VCC VCC u_muldiv.divisor\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_2532_ _0505_ _0503_ _0502_ VSS VSS VCC VCC _0507_ sky130_fd_sc_hd__nand3b_1
X_5251_ clknet_leaf_1_i_clk _0279_ VSS VSS VCC VCC u_muldiv.o_div\[28\] sky130_fd_sc_hd__dfxtp_2
X_2463_ net695 VSS VSS VCC VCC _0438_ sky130_fd_sc_hd__clkinv_2
X_4202_ net509 op_cnt\[0\] VSS VSS VCC VCC _0246_ sky130_fd_sc_hd__nor2_1
X_5182_ clknet_leaf_24_i_clk _0214_ VSS VSS VCC VCC u_muldiv.add_prev\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_4133_ _1831_ net378 net580 VSS VSS VCC VCC _1832_ sky130_fd_sc_hd__a21oi_1
X_4064_ net591 _1776_ _1777_ VSS VSS VCC VCC _1778_ sky130_fd_sc_hd__o21ba_1
X_3015_ net453 net611 _0812_ VSS VSS VCC VCC _0981_ sky130_fd_sc_hd__or3_1
X_4966_ _1138_ _1139_ net407 VSS VSS VCC VCC _0410_ sky130_fd_sc_hd__and3_2
X_3917_ u_pc_sel.i_pc_next\[8\] net122 net396 VSS VSS VCC VCC _0083_ sky130_fd_sc_hd__mux2_1
X_4897_ u_muldiv.divisor\[4\] net496 net342 u_muldiv.divisor\[5\] vssd1 vssd1 vccd1
+ vccd1 _0349_ sky130_fd_sc_hd__a22o_1
X_3848_ net508 _1667_ VSS VSS VCC VCC _1668_ sky130_fd_sc_hd__and2b_1
X_3779_ net502 net239 net723 _1617_ VSS VSS VCC VCC _0041_ sky130_fd_sc_hd__o211a_1
X_4820_ _2345_ u_muldiv.dividend\[25\] net433 VSS VSS VCC VCC _2362_ sky130_fd_sc_hd__a21oi_1
X_4751_ net684 net682 net679 _2267_ net371 VSS VSS VCC VCC _2299_ sky130_fd_sc_hd__o41a_1
X_3702_ net730 _1580_ net576 VSS VSS VCC VCC _1581_ sky130_fd_sc_hd__a21oi_4
X_4682_ _2234_ net372 net691 VSS VSS VCC VCC _2236_ sky130_fd_sc_hd__a21oi_1
X_3633_ net443 _1513_ _1516_ net733 VSS VSS VCC VCC _1517_ sky130_fd_sc_hd__a211o_2
X_3564_ net595 net697 net350 _1451_ VSS VSS VCC VCC _1452_ sky130_fd_sc_hd__o211ai_1
X_2515_ net641 net549 net678 net534 net424 VSS VSS VCC VCC _0490_ sky130_fd_sc_hd__o2111ai_2
X_5303_ clknet_4_8__leaf_i_clk _0331_ VSS VSS VCC VCC u_muldiv.dividend\[18\]
+ sky130_fd_sc_hd__dfxtp_4
X_3495_ net521 _1387_ net355 net210 VSS VSS VCC VCC _1388_ sky130_fd_sc_hd__a2bb2o_1
X_2446_ net616 VSS VSS VCC VCC _0421_ sky130_fd_sc_hd__inv_2
X_5234_ clknet_leaf_121_i_clk _0262_ VSS VSS VCC VCC u_muldiv.o_div\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_5165_ clknet_4_13__leaf_i_clk _0197_ VSS VSS VCC VCC u_muldiv.add_prev\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_4116_ net583 _1817_ _1818_ VSS VSS VCC VCC _1819_ sky130_fd_sc_hd__o21ba_1
X_5096_ clknet_leaf_177_i_clk _0129_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[11\]
+ sky130_fd_sc_hd__dfxtp_4
X_4047_ net596 net595 net594 _1753_ VSS VSS VCC VCC _1764_ sky130_fd_sc_hd__or4b_4
X_4949_ _1202_ _1203_ net407 VSS VSS VCC VCC _0393_ sky130_fd_sc_hd__and3_1
Xoutput280 net280 VSS VSS VCC VCC o_wdata[10] sky130_fd_sc_hd__buf_2
Xoutput291 net291 VSS VSS VCC VCC o_wdata[20] sky130_fd_sc_hd__buf_2
X_3280_ _0577_ _1212_ VSS VSS VCC VCC net194 sky130_fd_sc_hd__xor2_4
X_4803_ _2342_ u_muldiv.dividend\[24\] VSS VSS VCC VCC _2346_ sky130_fd_sc_hd__nand2_1
X_2995_ net661 u_muldiv.add_prev\[26\] net533 VSS VSS VCC VCC _0962_ sky130_fd_sc_hd__mux2_2
X_4734_ net462 _2262_ u_muldiv.dividend\[18\] VSS VSS VCC VCC _2283_ sky130_fd_sc_hd__o21ai_1
X_4665_ u_muldiv.dividend\[11\] _2220_ net318 VSS VSS VCC VCC _0324_ sky130_fd_sc_hd__mux2_1
X_3616_ u_muldiv.dividend\[13\] net420 net368 u_muldiv.o_div\[13\] net360 vssd1 vssd1
+ vccd1 vccd1 _1501_ sky130_fd_sc_hd__a221o_1
X_4596_ _2157_ _2156_ _2153_ _2154_ net439 VSS VSS VCC VCC _2158_ sky130_fd_sc_hd__o221a_1
X_3547_ net36 net731 net578 VSS VSS VCC VCC _1437_ sky130_fd_sc_hd__o21ba_1
X_3478_ net352 _1367_ _1368_ _1370_ net520 VSS VSS VCC VCC _1372_ sky130_fd_sc_hd__a41o_1
X_5217_ clknet_leaf_45_i_clk _0246_ VSS VSS VCC VCC op_cnt\[0\] sky130_fd_sc_hd__dfxtp_2
X_5148_ clknet_leaf_13_i_clk _0180_ VSS VSS VCC VCC u_muldiv.divisor\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_5079_ clknet_leaf_47_i_clk _0112_ VSS VSS VCC VCC u_muldiv.i_is_div sky130_fd_sc_hd__dfxtp_4
X_2780_ net568 net557 VSS VSS VCC VCC _0754_ sky130_fd_sc_hd__and2_1
X_4450_ _2058_ u_muldiv.o_div\[18\] VSS VSS VCC VCC _2061_ sky130_fd_sc_hd__nand2_1
X_3401_ net700 net697 net695 net694 net642 net627 VSS VSS VCC VCC _1298_ sky130_fd_sc_hd__mux4_1
X_4381_ u_muldiv.o_div\[2\] u_muldiv.o_div\[3\] u_muldiv.o_div\[4\] _1994_ vssd1 vssd1
+ vccd1 vccd1 _2006_ sky130_fd_sc_hd__or4_4
X_3332_ u_wr_mux.i_reg_data2\[8\] net279 net416 VSS VSS VCC VCC net309 sky130_fd_sc_hd__mux2_2
Xfanout709 u_bits.i_op1\[5\] VSS VSS VCC VCC net709 sky130_fd_sc_hd__clkbuf_4
X_3263_ _0660_ _1193_ _0681_ _0679_ _0738_ VSS VSS VCC VCC _1202_ sky130_fd_sc_hd__o221ai_4
X_5002_ clknet_leaf_11_i_clk _0035_ VSS VSS VCC VCC net277 sky130_fd_sc_hd__dfxtp_1
X_3194_ _0855_ _0850_ net616 VSS VSS VCC VCC _1150_ sky130_fd_sc_hd__mux2_1
X_2978_ net663 net664 net668 net670 net637 net625 VSS VSS VCC VCC _0946_ sky130_fd_sc_hd__mux4_1
X_4717_ _2267_ net373 net684 VSS VSS VCC VCC _2268_ sky130_fd_sc_hd__a21o_1
X_4648_ _1884_ _1887_ _2204_ VSS VSS VCC VCC _2205_ sky130_fd_sc_hd__a21oi_1
X_4579_ _1850_ _1851_ _1864_ _2141_ VSS VSS VCC VCC _2142_ sky130_fd_sc_hd__a31o_1
X_3950_ net530 net2 net394 VSS VSS VCC VCC _0113_ sky130_fd_sc_hd__mux2_1
X_2901_ net427 _0871_ VSS VSS VCC VCC _0872_ sky130_fd_sc_hd__xor2_1
X_3881_ net504 net93 net720 VSS VSS VCC VCC _1693_ sky130_fd_sc_hd__a21o_1
X_2832_ net609 net617 VSS VSS VCC VCC _0806_ sky130_fd_sc_hd__nor2_8
X_2763_ _0656_ _0659_ _0737_ VSS VSS VCC VCC _0738_ sky130_fd_sc_hd__o21ai_4
X_4502_ net316 _2099_ _2101_ VSS VSS VCC VCC _0280_ sky130_fd_sc_hd__a21oi_1
X_2694_ _0667_ _0668_ VSS VSS VCC VCC _0669_ sky130_fd_sc_hd__nand2_2
X_4433_ net436 _0455_ _2042_ net331 VSS VSS VCC VCC _2047_ sky130_fd_sc_hd__o31a_1
X_4364_ u_muldiv.outsign net483 _1989_ VSS VSS VCC VCC _1992_ sky130_fd_sc_hd__a21oi_4
Xfanout506 net507 VSS VSS VCC VCC net506 sky130_fd_sc_hd__buf_2
Xfanout517 net519 VSS VSS VCC VCC net517 sky130_fd_sc_hd__buf_8
X_3315_ _1236_ _1232_ _1244_ VSS VSS VCC VCC _1245_ sky130_fd_sc_hd__a21o_1
Xfanout528 net529 VSS VSS VCC VCC net528 sky130_fd_sc_hd__clkbuf_4
Xfanout539 net543 VSS VSS VCC VCC net539 sky130_fd_sc_hd__buf_6
X_4295_ _1911_ u_muldiv.dividend\[18\] VSS VSS VCC VCC _1923_ sky130_fd_sc_hd__nand2_1
X_3246_ _0638_ _0727_ _0733_ _0695_ VSS VSS VCC VCC _1189_ sky130_fd_sc_hd__a211o_1
X_3177_ net517 net523 _1132_ VSS VSS VCC VCC _1134_ sky130_fd_sc_hd__o21ai_1
X_3100_ net729 net26 _1061_ VSS VSS VCC VCC net265 sky130_fd_sc_hd__o21a_1
X_4080_ u_muldiv.divisor\[49\] net485 net336 u_muldiv.divisor\[50\] _1790_ vssd1 vssd1
+ vccd1 vccd1 _0169_ sky130_fd_sc_hd__a221o_1
X_3031_ _0993_ _0994_ _0995_ VSS VSS VCC VCC _0996_ sky130_fd_sc_hd__and3_1
Xinput180 i_reset_n VSS VSS VCC VCC net180 sky130_fd_sc_hd__buf_4
X_4982_ clknet_leaf_147_i_clk _0015_ VSS VSS VCC VCC u_bits.i_op1\[12\] sky130_fd_sc_hd__dfxtp_1
X_3933_ net228 net132 net390 VSS VSS VCC VCC _0096_ sky130_fd_sc_hd__mux2_1
X_3864_ net504 _1679_ VSS VSS VCC VCC _1680_ sky130_fd_sc_hd__and2b_1
X_2815_ net645 net713 VSS VSS VCC VCC _0789_ sky130_fd_sc_hd__nand2_1
X_3795_ net603 net624 net548 VSS VSS VCC VCC _1628_ sky130_fd_sc_hd__mux2_1
X_2746_ net449 net700 VSS VSS VCC VCC _0721_ sky130_fd_sc_hd__and2_1
X_2677_ net647 net552 net692 net542 net425 VSS VSS VCC VCC _0652_ sky130_fd_sc_hd__o2111ai_4
X_4416_ net322 _2031_ _2033_ u_muldiv.o_div\[11\] VSS VSS VCC VCC _0262_ sky130_fd_sc_hd__o22a_1
X_4347_ u_muldiv.divisor\[30\] _0447_ _1974_ VSS VSS VCC VCC _1975_ sky130_fd_sc_hd__o21a_1
Xfanout325 net326 VSS VSS VCC VCC net325 sky130_fd_sc_hd__buf_2
Xfanout336 net344 VSS VSS VCC VCC net336 sky130_fd_sc_hd__clkbuf_2
Xfanout347 _0890_ VSS VSS VCC VCC net347 sky130_fd_sc_hd__buf_4
Xfanout358 net359 VSS VSS VCC VCC net358 sky130_fd_sc_hd__clkbuf_4
Xfanout369 net370 VSS VSS VCC VCC net369 sky130_fd_sc_hd__clkbuf_4
X_4278_ _1902_ _1903_ _1904_ VSS VSS VCC VCC _1906_ sky130_fd_sc_hd__or3b_1
X_3229_ _0626_ _0631_ _0584_ _0603_ _0628_ VSS VSS VCC VCC _1176_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_139_i_clk clknet_4_10__leaf_i_clk VSS VSS VCC VCC clknet_leaf_139_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2600_ net449 net460 VSS VSS VCC VCC _0575_ sky130_fd_sc_hd__and2_1
X_3580_ _1006_ net603 VSS VSS VCC VCC _1467_ sky130_fd_sc_hd__nand2b_1
X_2531_ _0504_ _0505_ VSS VSS VCC VCC _0506_ sky130_fd_sc_hd__nand2_1
X_5250_ clknet_leaf_2_i_clk _0278_ VSS VSS VCC VCC u_muldiv.o_div\[27\] sky130_fd_sc_hd__dfxtp_1
X_2462_ net697 VSS VSS VCC VCC _0437_ sky130_fd_sc_hd__clkinv_2
X_4201_ net183 u_muldiv.mul\[30\] net405 VSS VSS VCC VCC _0245_ sky130_fd_sc_hd__mux2_1
X_5181_ clknet_leaf_58_i_clk _0213_ VSS VSS VCC VCC u_muldiv.add_prev\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_56_i_clk clknet_4_6__leaf_i_clk VSS VSS VCC VCC clknet_leaf_56_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4132_ u_bits.i_op2\[28\] net581 _1823_ VSS VSS VCC VCC _1831_ sky130_fd_sc_hd__or3_1
X_4063_ _1775_ net381 net591 net330 VSS VSS VCC VCC _1777_ sky130_fd_sc_hd__a31o_1
X_3014_ _0804_ _0810_ net453 VSS VSS VCC VCC _0980_ sky130_fd_sc_hd__mux2_1
X_4965_ net549 net499 _1109_ _1110_ VSS VSS VCC VCC _0409_ sky130_fd_sc_hd__nor4_1
X_3916_ u_pc_sel.i_pc_next\[7\] net121 net394 VSS VSS VCC VCC _0082_ sky130_fd_sc_hd__mux2_1
X_4896_ u_muldiv.divisor\[3\] net497 net343 u_muldiv.divisor\[4\] vssd1 vssd1 vccd1
+ vccd1 _0348_ sky130_fd_sc_hd__a22o_1
X_3847_ net589 net591 net547 VSS VSS VCC VCC _1667_ sky130_fd_sc_hd__mux2_1
X_3778_ net143 net511 VSS VSS VCC VCC _1617_ sky130_fd_sc_hd__nand2b_1
X_2729_ _0698_ _0699_ _0701_ VSS VSS VCC VCC _0704_ sky130_fd_sc_hd__a21oi_1
X_5379_ clknet_leaf_156_i_clk _0406_ VSS VSS VCC VCC u_muldiv.mul\[58\] sky130_fd_sc_hd__dfxtp_1
X_4750_ u_muldiv.dividend\[19\] _2284_ VSS VSS VCC VCC _2298_ sky130_fd_sc_hd__nor2_1
X_3701_ net527 _1571_ _1579_ VSS VSS VCC VCC _1580_ sky130_fd_sc_hd__a21o_1
X_4681_ _2234_ net372 net690 VSS VSS VCC VCC _2235_ sky130_fd_sc_hd__and3_1
X_3632_ net556 u_muldiv.mul\[14\] net415 net528 _1515_ VSS VSS VCC VCC _1516_
+ sky130_fd_sc_hd__o311a_1
X_3563_ net566 _0437_ net595 VSS VSS VCC VCC _1451_ sky130_fd_sc_hd__or3b_1
X_5302_ clknet_4_8__leaf_i_clk _0330_ VSS VSS VCC VCC u_muldiv.dividend\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_2514_ _0480_ _0488_ _0481_ VSS VSS VCC VCC _0489_ sky130_fd_sc_hd__a21bo_1
X_3494_ net353 _1382_ _1383_ _1385_ _1386_ VSS VSS VCC VCC _1387_ sky130_fd_sc_hd__a41o_1
X_5233_ clknet_leaf_121_i_clk _0261_ VSS VSS VCC VCC u_muldiv.o_div\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_2445_ net620 VSS VSS VCC VCC _0420_ sky130_fd_sc_hd__clkinv_2
X_5164_ clknet_leaf_74_i_clk _0196_ VSS VSS VCC VCC u_muldiv.add_prev\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4115_ _1816_ net382 net583 net329 VSS VSS VCC VCC _1818_ sky130_fd_sc_hd__a31o_1
X_5095_ clknet_leaf_60_i_clk _0128_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_4046_ u_muldiv.divisor\[42\] net484 net335 net737 _1763_ VSS VSS VCC VCC
+ _0162_ sky130_fd_sc_hd__a221o_1
X_4948_ _1194_ _1195_ net406 VSS VSS VCC VCC _0392_ sky130_fd_sc_hd__and3_1
X_4879_ net652 _2415_ net383 VSS VSS VCC VCC _2416_ sky130_fd_sc_hd__o21ai_1
Xoutput270 net270 VSS VSS VCC VCC o_result[3] sky130_fd_sc_hd__buf_2
Xoutput281 net281 VSS VSS VCC VCC o_wdata[11] sky130_fd_sc_hd__buf_2
Xoutput292 net292 VSS VSS VCC VCC o_wdata[21] sky130_fd_sc_hd__buf_2
X_4802_ u_muldiv.dividend\[24\] u_muldiv.dividend\[23\] u_muldiv.dividend\[22\] _2322_
+ VSS VSS VCC VCC _2345_ sky130_fd_sc_hd__or4_4
X_2994_ net516 net523 _0959_ VSS VSS VCC VCC _0961_ sky130_fd_sc_hd__o21ai_2
X_4733_ u_muldiv.dividend\[17\] net319 _2282_ VSS VSS VCC VCC _0330_ sky130_fd_sc_hd__o21a_1
X_4664_ net437 _2214_ _2217_ _2218_ _2219_ VSS VSS VCC VCC _2220_ sky130_fd_sc_hd__a32o_1
X_3615_ net521 _1498_ _1499_ net356 _1196_ VSS VSS VCC VCC _1500_ sky130_fd_sc_hd__o32a_1
X_4595_ net709 _2155_ net459 VSS VSS VCC VCC _2157_ sky130_fd_sc_hd__o21ai_1
X_3546_ net443 _1432_ _1435_ net734 VSS VSS VCC VCC _1436_ sky130_fd_sc_hd__a211o_1
X_3477_ net607 net710 net352 VSS VSS VCC VCC _1371_ sky130_fd_sc_hd__a21oi_1
X_5216_ clknet_leaf_40_i_clk _0000_ VSS VSS VCC VCC u_muldiv.i_on_end sky130_fd_sc_hd__dfxtp_4
X_5147_ clknet_leaf_12_i_clk _0179_ VSS VSS VCC VCC u_muldiv.divisor\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_5078_ clknet_leaf_116_i_clk _0111_ VSS VSS VCC VCC net217 sky130_fd_sc_hd__dfxtp_1
X_4029_ net599 net598 _1741_ net379 VSS VSS VCC VCC _1750_ sky130_fd_sc_hd__o31a_1
X_3400_ net690 net688 net686 net684 net642 net627 VSS VSS VCC VCC _1297_ sky130_fd_sc_hd__mux4_2
X_4380_ u_muldiv.o_div\[0\] u_muldiv.o_div\[1\] u_muldiv.o_div\[2\] u_muldiv.o_div\[3\]
+ VSS VSS VCC VCC _2005_ sky130_fd_sc_hd__or4_1
X_3331_ _1248_ net400 _1257_ VSS VSS VCC VCC _0003_ sky130_fd_sc_hd__a21oi_1
X_3262_ _1201_ VSS VSS VCC VCC net189 sky130_fd_sc_hd__inv_4
X_5001_ clknet_leaf_11_i_clk _0034_ VSS VSS VCC VCC u_bits.i_op1\[31\] sky130_fd_sc_hd__dfxtp_2
X_3193_ net328 _0842_ net347 _1148_ net411 VSS VSS VCC VCC _1149_ sky130_fd_sc_hd__a311o_1
X_2977_ net620 _0944_ _0943_ VSS VSS VCC VCC _0945_ sky130_fd_sc_hd__o21ai_4
X_4716_ net690 net688 net686 _2234_ VSS VSS VCC VCC _2267_ sky130_fd_sc_hd__or4_2
X_4647_ _1884_ _1887_ net471 VSS VSS VCC VCC _2204_ sky130_fd_sc_hd__o21ai_1
X_4578_ _2140_ net473 VSS VSS VCC VCC _2141_ sky130_fd_sc_hd__nand2_1
X_3529_ u_muldiv.o_div\[7\] net366 net358 _1419_ VSS VSS VCC VCC _1420_ sky130_fd_sc_hd__a211o_1
X_2900_ net445 u_bits.i_op2\[24\] _0464_ net666 VSS VSS VCC VCC _0871_ sky130_fd_sc_hd__a22o_1
X_3880_ net504 _1691_ VSS VSS VCC VCC _1692_ sky130_fd_sc_hd__and2b_1
X_2831_ _0803_ _0801_ _0800_ _0798_ net630 net621 VSS VSS VCC VCC _0805_ sky130_fd_sc_hd__mux4_2
X_2762_ _0646_ _0658_ VSS VSS VCC VCC _0737_ sky130_fd_sc_hd__nand2_1
X_4501_ net316 _2100_ u_muldiv.o_div\[29\] VSS VSS VCC VCC _2101_ sky130_fd_sc_hd__a21oi_1
X_2693_ net687 u_muldiv.add_prev\[15\] net542 VSS VSS VCC VCC _0668_ sky130_fd_sc_hd__mux2_1
X_4432_ u_muldiv.o_div\[14\] net318 _2046_ VSS VSS VCC VCC _0265_ sky130_fd_sc_hd__o21a_1
X_4363_ u_muldiv.outsign net483 VSS VSS VCC VCC _1991_ sky130_fd_sc_hd__nand2_8
Xfanout507 net508 VSS VSS VCC VCC net507 sky130_fd_sc_hd__buf_2
Xfanout518 net519 VSS VSS VCC VCC net518 sky130_fd_sc_hd__buf_6
X_3314_ _1240_ _1243_ net561 VSS VSS VCC VCC _1244_ sky130_fd_sc_hd__o21bai_1
Xfanout529 net530 VSS VSS VCC VCC net529 sky130_fd_sc_hd__clkbuf_4
X_4294_ _1916_ _1921_ _1909_ _1912_ VSS VSS VCC VCC _1922_ sky130_fd_sc_hd__a211o_1
X_3245_ _1188_ VSS VSS VCC VCC net185 sky130_fd_sc_hd__inv_2
X_3176_ net517 net523 _1132_ VSS VSS VCC VCC _1133_ sky130_fd_sc_hd__or3_1
X_3030_ net659 u_muldiv.add_prev\[27\] net533 VSS VSS VCC VCC _0995_ sky130_fd_sc_hd__mux2_1
Xinput170 i_reg_data2[4] VSS VSS VCC VCC net170 sky130_fd_sc_hd__clkbuf_1
Xinput181 i_store VSS VSS VCC VCC net181 sky130_fd_sc_hd__clkbuf_1
X_4981_ clknet_leaf_134_i_clk _0014_ VSS VSS VCC VCC u_bits.i_op1\[11\] sky130_fd_sc_hd__dfxtp_4
X_3932_ net227 net131 net393 VSS VSS VCC VCC _0095_ sky130_fd_sc_hd__mux2_1
X_3863_ u_bits.i_op2\[21\] net587 net546 VSS VSS VCC VCC _1679_ sky130_fd_sc_hd__mux2_1
X_2814_ _0419_ net706 _0787_ VSS VSS VCC VCC _0788_ sky130_fd_sc_hd__a21oi_1
X_3794_ net624 net724 _1627_ _1626_ VSS VSS VCC VCC _0046_ sky130_fd_sc_hd__o22a_1
X_2745_ net541 u_muldiv.add_prev\[9\] VSS VSS VCC VCC _0720_ sky130_fd_sc_hd__and2_1
X_2676_ net542 net692 VSS VSS VCC VCC _0651_ sky130_fd_sc_hd__and2_1
X_4415_ net324 net375 _2028_ _2032_ VSS VSS VCC VCC _2033_ sky130_fd_sc_hd__o2bb2a_1
X_4346_ u_muldiv.divisor\[31\] u_muldiv.dividend\[31\] VSS VSS VCC VCC _1974_
+ sky130_fd_sc_hd__nand2b_1
Xfanout315 net317 VSS VSS VCC VCC net315 sky130_fd_sc_hd__clkbuf_8
Xfanout326 _1990_ VSS VSS VCC VCC net326 sky130_fd_sc_hd__buf_6
Xfanout337 net344 VSS VSS VCC VCC net337 sky130_fd_sc_hd__clkbuf_4
Xfanout348 _0785_ VSS VSS VCC VCC net348 sky130_fd_sc_hd__clkbuf_8
Xfanout359 net360 VSS VSS VCC VCC net359 sky130_fd_sc_hd__clkbuf_4
X_4277_ _1903_ _1904_ VSS VSS VCC VCC _1905_ sky130_fd_sc_hd__nand2b_1
X_3228_ _1175_ VSS VSS VCC VCC net212 sky130_fd_sc_hd__clkinv_2
X_3159_ net601 _1113_ _1116_ VSS VSS VCC VCC _1117_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_4_6__f_i_clk clknet_2_1_0_i_clk VSS VSS VCC VCC clknet_4_6__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2530_ net681 u_muldiv.add_prev\[18\] net536 VSS VSS VCC VCC _0505_ sky130_fd_sc_hd__mux2_1
X_2461_ net704 VSS VSS VCC VCC _0436_ sky130_fd_sc_hd__inv_2
X_4200_ u_muldiv.mul\[30\] u_muldiv.mul\[29\] net405 VSS VSS VCC VCC _0244_
+ sky130_fd_sc_hd__mux2_1
X_5180_ clknet_leaf_56_i_clk _0212_ VSS VSS VCC VCC u_muldiv.add_prev\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_4131_ u_muldiv.divisor\[60\] net482 net337 u_muldiv.divisor\[61\] _1830_ vssd1 vssd1
+ vccd1 vccd1 _0180_ sky130_fd_sc_hd__a221o_1
X_4062_ _1774_ u_bits.i_op2\[12\] _1764_ net381 VSS VSS VCC VCC _1776_ sky130_fd_sc_hd__o31a_1
X_3013_ _0897_ _0794_ net613 _0978_ VSS VSS VCC VCC _0979_ sky130_fd_sc_hd__o22a_2
X_4964_ _1071_ _1072_ net407 VSS VSS VCC VCC _0408_ sky130_fd_sc_hd__and3_2
X_3915_ u_pc_sel.i_pc_next\[6\] net120 net397 VSS VSS VCC VCC _0081_ sky130_fd_sc_hd__mux2_1
X_4895_ u_muldiv.divisor\[2\] net498 net343 u_muldiv.divisor\[3\] vssd1 vssd1 vccd1
+ vccd1 _0347_ sky130_fd_sc_hd__a22o_1
X_3846_ net591 net727 _1666_ _1665_ VSS VSS VCC VCC _0059_ sky130_fd_sc_hd__o22a_1
X_3777_ net509 net238 net727 _1616_ VSS VSS VCC VCC _0040_ sky130_fd_sc_hd__o211a_1
X_2728_ net428 _0696_ _0697_ _0701_ VSS VSS VCC VCC _0703_ sky130_fd_sc_hd__a31o_1
X_2659_ _0614_ _0615_ _0626_ _0631_ VSS VSS VCC VCC _0634_ sky130_fd_sc_hd__and4_2
X_5378_ clknet_leaf_156_i_clk _0405_ VSS VSS VCC VCC u_muldiv.mul\[57\] sky130_fd_sc_hd__dfxtp_1
X_4329_ u_muldiv.divisor\[25\] _0449_ _1956_ VSS VSS VCC VCC _1957_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_170_i_clk clknet_4_0__leaf_i_clk VSS VSS VCC VCC clknet_leaf_170_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout690 net691 VSS VSS VCC VCC net690 sky130_fd_sc_hd__buf_4
X_3700_ net521 _1578_ net356 _1208_ net446 VSS VSS VCC VCC _1579_ sky130_fd_sc_hd__o221a_2
X_4680_ _2206_ _0439_ _0438_ _0437_ VSS VSS VCC VCC _2234_ sky130_fd_sc_hd__nand4_4
X_3631_ u_muldiv.o_div\[14\] net366 net358 _1514_ VSS VSS VCC VCC _1515_ sky130_fd_sc_hd__a211o_1
X_3562_ _1450_ u_pc_sel.i_pc_next\[9\] net577 VSS VSS VCC VCC net276 sky130_fd_sc_hd__mux2_2
X_5301_ clknet_4_8__leaf_i_clk _0329_ VSS VSS VCC VCC u_muldiv.dividend\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_2513_ _0484_ _0485_ _0487_ VSS VSS VCC VCC _0488_ sky130_fd_sc_hd__a21o_2
X_3493_ u_bits.i_op2\[5\] net709 net353 VSS VSS VCC VCC _1386_ sky130_fd_sc_hd__a21oi_1
X_5232_ clknet_leaf_121_i_clk _0260_ VSS VSS VCC VCC u_muldiv.o_div\[9\] sky130_fd_sc_hd__dfxtp_2
X_2444_ net645 VSS VSS VCC VCC _0419_ sky130_fd_sc_hd__inv_4
X_5163_ clknet_leaf_74_i_clk _0195_ VSS VSS VCC VCC u_muldiv.add_prev\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4114_ net586 net585 net584 _1806_ net378 VSS VSS VCC VCC _1817_ sky130_fd_sc_hd__o41a_1
X_5094_ clknet_leaf_132_i_clk _0127_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[9\]
+ sky130_fd_sc_hd__dfxtp_4
X_4045_ _1761_ _1762_ VSS VSS VCC VCC _1763_ sky130_fd_sc_hd__nor2_1
X_4947_ _1193_ _1197_ net406 VSS VSS VCC VCC _0391_ sky130_fd_sc_hd__and3_1
X_4878_ net654 _2404_ net370 VSS VSS VCC VCC _2415_ sky130_fd_sc_hd__o21ai_1
X_3829_ net505 net79 net719 VSS VSS VCC VCC _1654_ sky130_fd_sc_hd__a21o_1
Xoutput260 net260 VSS VSS VCC VCC o_result[23] sky130_fd_sc_hd__buf_2
Xoutput271 net271 VSS VSS VCC VCC o_result[4] sky130_fd_sc_hd__buf_2
Xoutput282 net282 VSS VSS VCC VCC o_wdata[12] sky130_fd_sc_hd__buf_2
Xoutput293 net293 VSS VSS VCC VCC o_wdata[22] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_40_i_clk clknet_4_5__leaf_i_clk VSS VSS VCC VCC clknet_leaf_40_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_2_0_0_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_55_i_clk clknet_4_7__leaf_i_clk VSS VSS VCC VCC clknet_leaf_55_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4801_ u_muldiv.dividend\[23\] _2344_ net317 VSS VSS VCC VCC _0336_ sky130_fd_sc_hd__mux2_1
X_2993_ net533 net661 _0463_ _0958_ net427 VSS VSS VCC VCC _0960_ sky130_fd_sc_hd__a311o_2
X_4732_ _2281_ _2280_ _2279_ net319 VSS VSS VCC VCC _2282_ sky130_fd_sc_hd__o211ai_1
X_4663_ _2201_ u_muldiv.dividend\[11\] net435 VSS VSS VCC VCC _2219_ sky130_fd_sc_hd__a21oi_1
X_3614_ u_bits.i_op2\[13\] net691 net352 VSS VSS VCC VCC _1499_ sky130_fd_sc_hd__a21oi_1
X_4594_ net712 u_bits.i_op1\[4\] _2131_ net374 net709 VSS VSS VCC VCC _2156_
+ sky130_fd_sc_hd__o311a_1
X_3545_ net559 u_muldiv.mul\[8\] net413 net528 _1434_ VSS VSS VCC VCC _1435_
+ sky130_fd_sc_hd__o311a_1
X_3476_ net607 net710 net350 _1369_ VSS VSS VCC VCC _1370_ sky130_fd_sc_hd__o211ai_1
X_5215_ clknet_leaf_58_i_clk _0002_ VSS VSS VCC VCC u_muldiv.i_on_wait sky130_fd_sc_hd__dfxtp_2
X_5146_ clknet_leaf_29_i_clk _0178_ VSS VSS VCC VCC u_muldiv.divisor\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_5077_ clknet_leaf_10_i_clk _0110_ VSS VSS VCC VCC net216 sky130_fd_sc_hd__dfxtp_4
X_4028_ net600 net599 net598 _1737_ VSS VSS VCC VCC _1749_ sky130_fd_sc_hd__or4_1
X_3330_ net40 net41 net407 VSS VSS VCC VCC _1257_ sky130_fd_sc_hd__and3_1
X_3261_ _0671_ _1200_ VSS VSS VCC VCC _1201_ sky130_fd_sc_hd__xnor2_4
X_5000_ clknet_leaf_84_i_clk _0033_ VSS VSS VCC VCC u_bits.i_op1\[30\] sky130_fd_sc_hd__dfxtp_1
X_3192_ net561 _1146_ _1147_ net349 VSS VSS VCC VCC _1148_ sky130_fd_sc_hd__o211a_1
X_2976_ net682 net684 net686 net688 net642 net631 VSS VSS VCC VCC _0944_ sky130_fd_sc_hd__mux4_2
X_4715_ net690 net688 net686 _2234_ VSS VSS VCC VCC _2266_ sky130_fd_sc_hd__nor4_1
X_4646_ _1884_ _1887_ VSS VSS VCC VCC _2203_ sky130_fd_sc_hd__nor2_1
X_4577_ _1850_ _1851_ _1864_ VSS VSS VCC VCC _2140_ sky130_fd_sc_hd__a21o_1
X_3528_ net566 net556 u_muldiv.dividend\[7\] u_muldiv.mul\[39\] net362 vssd1 vssd1
+ vccd1 vccd1 _1419_ sky130_fd_sc_hd__a32o_1
X_3459_ net441 u_muldiv.mul\[35\] net414 _1353_ VSS VSS VCC VCC _1354_ sky130_fd_sc_hd__a31o_1
X_5129_ clknet_leaf_37_i_clk _0161_ VSS VSS VCC VCC u_muldiv.divisor\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_2830_ net689 net690 net693 net695 net642 net627 VSS VSS VCC VCC _0804_ sky130_fd_sc_hd__mux4_1
X_2761_ _0706_ _0734_ _0735_ VSS VSS VCC VCC _0736_ sky130_fd_sc_hd__o21ai_4
X_4500_ _2095_ u_muldiv.quotient_msk\[29\] net434 VSS VSS VCC VCC _2100_ sky130_fd_sc_hd__mux2_1
X_2692_ _0665_ _0666_ VSS VSS VCC VCC _0667_ sky130_fd_sc_hd__nand2_1
X_4431_ _2043_ _2044_ _2045_ net319 VSS VSS VCC VCC _2046_ sky130_fd_sc_hd__o211ai_1
X_4362_ _1973_ _1975_ net466 _1988_ VSS VSS VCC VCC _1990_ sky130_fd_sc_hd__a31o_4
X_3313_ _1238_ _1241_ net440 VSS VSS VCC VCC _1243_ sky130_fd_sc_hd__a21o_1
Xfanout508 net240 VSS VSS VCC VCC net508 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout519 u_muldiv.i_op2_signed VSS VSS VCC VCC net519 sky130_fd_sc_hd__clkbuf_8
X_4293_ u_muldiv.divisor\[16\] _1917_ u_muldiv.dividend\[16\] VSS VSS VCC VCC
+ _1921_ sky130_fd_sc_hd__or3b_1
X_3244_ _1186_ _1187_ VSS VSS VCC VCC _1188_ sky130_fd_sc_hd__nand2_4
X_3175_ net532 u_bits.i_op2\[31\] _1131_ VSS VSS VCC VCC _1132_ sky130_fd_sc_hd__o21ai_2
X_2959_ _0920_ _0927_ VSS VSS VCC VCC _0928_ sky130_fd_sc_hd__xnor2_4
X_4629_ _1879_ _2183_ net471 net494 VSS VSS VCC VCC _2188_ sky130_fd_sc_hd__a31o_1
Xinput160 i_reg_data2[24] VSS VSS VCC VCC net160 sky130_fd_sc_hd__buf_2
Xinput171 i_reg_data2[5] VSS VSS VCC VCC net171 sky130_fd_sc_hd__clkbuf_1
Xinput182 i_to_trap VSS VSS VCC VCC net182 sky130_fd_sc_hd__clkbuf_4
X_4980_ clknet_leaf_74_i_clk _0013_ VSS VSS VCC VCC u_bits.i_op1\[10\] sky130_fd_sc_hd__dfxtp_1
X_3931_ net226 net130 net388 VSS VSS VCC VCC _0094_ sky130_fd_sc_hd__mux2_1
X_3862_ net587 net728 _1678_ _1677_ VSS VSS VCC VCC _0063_ sky130_fd_sc_hd__o22a_1
X_2813_ net645 net708 VSS VSS VCC VCC _0787_ sky130_fd_sc_hd__and2_1
X_3793_ net501 net99 net720 VSS VSS VCC VCC _1627_ sky130_fd_sc_hd__a21o_1
X_2744_ net518 net526 _0717_ VSS VSS VCC VCC _0719_ sky130_fd_sc_hd__o21ai_2
X_2675_ _0649_ VSS VSS VCC VCC _0650_ sky130_fd_sc_hd__inv_2
X_4414_ net435 u_muldiv.quotient_msk\[11\] VSS VSS VCC VCC _2032_ sky130_fd_sc_hd__and2_1
X_4345_ _1970_ _1971_ _1969_ VSS VSS VCC VCC _1973_ sky130_fd_sc_hd__o21ai_4
Xfanout316 net317 VSS VSS VCC VCC net316 sky130_fd_sc_hd__clkbuf_2
Xfanout327 _0769_ VSS VSS VCC VCC net327 sky130_fd_sc_hd__buf_4
Xfanout338 net340 VSS VSS VCC VCC net338 sky130_fd_sc_hd__buf_4
Xfanout349 _0785_ VSS VSS VCC VCC net349 sky130_fd_sc_hd__clkbuf_4
X_4276_ u_muldiv.dividend\[15\] u_muldiv.divisor\[15\] VSS VSS VCC VCC _1904_
+ sky130_fd_sc_hd__nand2b_1
X_3227_ _1173_ _1174_ VSS VSS VCC VCC _1175_ sky130_fd_sc_hd__nand2_4
X_3158_ net601 _1115_ _0814_ VSS VSS VCC VCC _1116_ sky130_fd_sc_hd__o21ai_1
X_3089_ _0905_ _0906_ net346 _1050_ net345 VSS VSS VCC VCC _1051_ sky130_fd_sc_hd__o221ai_1
X_2460_ net710 VSS VSS VCC VCC _0435_ sky130_fd_sc_hd__inv_2
X_4130_ _1828_ _1829_ VSS VSS VCC VCC _1830_ sky130_fd_sc_hd__nor2_1
X_4061_ net594 _1774_ u_bits.i_op2\[12\] _1760_ VSS VSS VCC VCC _1775_ sky130_fd_sc_hd__or4_1
X_3012_ _0788_ _0790_ _0800_ _0798_ net629 net454 VSS VSS VCC VCC _0978_ sky130_fd_sc_hd__mux4_1
X_4963_ net547 net203 _0432_ VSS VSS VCC VCC _0407_ sky130_fd_sc_hd__and3b_1
X_3914_ u_pc_sel.i_pc_next\[5\] net119 net387 VSS VSS VCC VCC _0080_ sky130_fd_sc_hd__mux2_1
X_4894_ u_muldiv.divisor\[1\] net498 net343 u_muldiv.divisor\[2\] vssd1 vssd1 vccd1
+ vccd1 _0346_ sky130_fd_sc_hd__a22o_1
X_3845_ net512 net83 net722 VSS VSS VCC VCC _1666_ sky130_fd_sc_hd__a21o_1
X_3776_ net142 net509 VSS VSS VCC VCC _1616_ sky130_fd_sc_hd__nand2b_1
X_2727_ _0698_ _0699_ _0701_ VSS VSS VCC VCC _0702_ sky130_fd_sc_hd__nand3_2
X_2658_ _0626_ _0631_ VSS VSS VCC VCC _0633_ sky130_fd_sc_hd__nand2_1
X_2589_ net447 net634 VSS VSS VCC VCC _0564_ sky130_fd_sc_hd__nand2_1
X_5377_ clknet_leaf_157_i_clk _0404_ VSS VSS VCC VCC u_muldiv.mul\[56\] sky130_fd_sc_hd__dfxtp_1
X_4328_ u_muldiv.divisor\[25\] _0449_ _1945_ VSS VSS VCC VCC _1956_ sky130_fd_sc_hd__a21oi_1
X_4259_ _1885_ _1886_ VSS VSS VCC VCC _1887_ sky130_fd_sc_hd__or2_1
Xfanout680 net681 VSS VSS VCC VCC net680 sky130_fd_sc_hd__buf_4
Xfanout691 net692 VSS VSS VCC VCC net691 sky130_fd_sc_hd__buf_4
X_3630_ net567 net556 u_muldiv.dividend\[14\] u_muldiv.mul\[46\] net362 vssd1 vssd1
+ vccd1 vccd1 _1514_ sky130_fd_sc_hd__a32o_1
X_3561_ _1449_ net37 net734 VSS VSS VCC VCC _1450_ sky130_fd_sc_hd__mux2_1
X_5300_ clknet_leaf_143_i_clk _0328_ VSS VSS VCC VCC u_muldiv.dividend\[15\]
+ sky130_fd_sc_hd__dfxtp_4
X_2512_ net446 net676 _0486_ VSS VSS VCC VCC _0487_ sky130_fd_sc_hd__a21oi_1
X_3492_ net600 net709 net351 _1384_ VSS VSS VCC VCC _1385_ sky130_fd_sc_hd__o211ai_1
X_2443_ u_muldiv.divisor\[1\] VSS VSS VCC VCC _0418_ sky130_fd_sc_hd__inv_2
X_5231_ clknet_leaf_118_i_clk _0259_ VSS VSS VCC VCC u_muldiv.o_div\[8\] sky130_fd_sc_hd__dfxtp_2
X_5162_ clknet_leaf_77_i_clk _0194_ VSS VSS VCC VCC u_muldiv.add_prev\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4113_ net586 net585 net584 _1806_ VSS VSS VCC VCC _1816_ sky130_fd_sc_hd__or4_2
X_5093_ clknet_leaf_83_i_clk _0126_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[8\]
+ sky130_fd_sc_hd__dfxtp_4
X_4044_ _1760_ net381 net594 net330 VSS VSS VCC VCC _1762_ sky130_fd_sc_hd__a31o_1
X_4946_ _1186_ _1187_ net407 VSS VSS VCC VCC _0390_ sky130_fd_sc_hd__and3_1
X_4877_ _2412_ _2413_ net479 VSS VSS VCC VCC _2414_ sky130_fd_sc_hd__o21ai_1
X_3828_ net505 _1652_ VSS VSS VCC VCC _1653_ sky130_fd_sc_hd__and2b_1
X_3759_ net662 net62 net388 VSS VSS VCC VCC _0028_ sky130_fd_sc_hd__mux2_1
Xoutput250 net250 VSS VSS VCC VCC o_result[14] sky130_fd_sc_hd__buf_2
Xoutput261 net261 VSS VSS VCC VCC o_result[24] sky130_fd_sc_hd__buf_2
Xoutput272 net272 VSS VSS VCC VCC o_result[5] sky130_fd_sc_hd__buf_2
Xoutput283 net283 VSS VSS VCC VCC o_wdata[13] sky130_fd_sc_hd__buf_2
Xoutput294 net294 VSS VSS VCC VCC o_wdata[23] sky130_fd_sc_hd__buf_2
X_4800_ net480 _2342_ _2343_ _2337_ _2341_ VSS VSS VCC VCC _2344_ sky130_fd_sc_hd__a32o_1
X_2992_ net533 net661 _0463_ _0958_ VSS VSS VCC VCC _0959_ sky130_fd_sc_hd__a31o_1
X_4731_ _2262_ net462 net437 VSS VSS VCC VCC _2281_ sky130_fd_sc_hd__a21o_1
X_4662_ u_muldiv.dividend\[11\] u_muldiv.dividend\[10\] u_muldiv.dividend\[9\] _2180_
+ VSS VSS VCC VCC _2218_ sky130_fd_sc_hd__or4_1
X_3613_ _1494_ _1496_ _1497_ VSS VSS VCC VCC _1498_ sky130_fd_sc_hd__a21oi_2
X_4593_ net713 net711 _2131_ net374 VSS VSS VCC VCC _2155_ sky130_fd_sc_hd__o31a_1
X_3544_ u_muldiv.o_div\[8\] net366 net358 _1433_ VSS VSS VCC VCC _1434_ sky130_fd_sc_hd__a211o_1
X_3475_ net566 _0435_ net607 VSS VSS VCC VCC _1369_ sky130_fd_sc_hd__or3b_1
X_5214_ clknet_leaf_55_i_clk _0001_ VSS VSS VCC VCC net240 sky130_fd_sc_hd__dfxtp_4
X_5145_ clknet_leaf_29_i_clk _0177_ VSS VSS VCC VCC u_muldiv.divisor\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_5076_ clknet_leaf_9_i_clk _0109_ VSS VSS VCC VCC net215 sky130_fd_sc_hd__dfxtp_4
X_4027_ u_muldiv.divisor\[38\] net482 net337 u_muldiv.divisor\[39\] _1748_ vssd1 vssd1
+ vccd1 vccd1 _0158_ sky130_fd_sc_hd__a221o_1
X_4929_ u_muldiv.quotient_msk\[0\] _1989_ u_muldiv.o_div\[0\] VSS VSS VCC VCC
+ _2432_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_122_i_clk clknet_4_11__leaf_i_clk VSS VSS VCC VCC clknet_leaf_122_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_137_i_clk clknet_4_8__leaf_i_clk VSS VSS VCC VCC clknet_leaf_137_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3260_ _0680_ _0738_ _1199_ _0681_ VSS VSS VCC VCC _1200_ sky130_fd_sc_hd__a31o_1
X_3191_ net651 u_bits.i_op2\[31\] VSS VSS VCC VCC _1147_ sky130_fd_sc_hd__or2_1
X_2975_ net454 _0942_ VSS VSS VCC VCC _0943_ sky130_fd_sc_hd__or2_1
X_4714_ _1908_ _1915_ _2264_ VSS VSS VCC VCC _2265_ sky130_fd_sc_hd__o21a_1
X_4645_ _2200_ _2201_ net435 VSS VSS VCC VCC _2202_ sky130_fd_sc_hd__a21o_1
X_4576_ u_muldiv.dividend\[3\] _2139_ net320 VSS VSS VCC VCC _0316_ sky130_fd_sc_hd__mux2_1
X_3527_ net520 _1416_ _1417_ net356 _1175_ VSS VSS VCC VCC _1418_ sky130_fd_sc_hd__o32ai_4
X_3458_ u_muldiv.dividend\[3\] net421 net367 u_muldiv.o_div\[3\] net358 vssd1 vssd1
+ vccd1 vccd1 _1353_ sky130_fd_sc_hd__a221o_1
X_3389_ _1269_ _1285_ _1286_ VSS VSS VCC VCC _1287_ sky130_fd_sc_hd__a21oi_2
X_5128_ clknet_leaf_37_i_clk _0160_ VSS VSS VCC VCC u_muldiv.divisor\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_5059_ clknet_leaf_116_i_clk _0092_ VSS VSS VCC VCC net243 sky130_fd_sc_hd__dfxtp_4
X_2760_ _0693_ _0704_ _0702_ VSS VSS VCC VCC _0735_ sky130_fd_sc_hd__o21a_1
X_2691_ net519 net526 _0663_ _0664_ VSS VSS VCC VCC _0666_ sky130_fd_sc_hd__o211ai_2
X_4430_ u_muldiv.quotient_msk\[14\] u_muldiv.o_div\[14\] net340 vssd1 vssd1 vccd1
+ vccd1 _2045_ sky130_fd_sc_hd__o21ai_1
X_4361_ _1973_ _1975_ net466 _1988_ VSS VSS VCC VCC _1989_ sky130_fd_sc_hd__a31oi_4
X_3312_ _1238_ _1241_ VSS VSS VCC VCC _1242_ sky130_fd_sc_hd__nand2_1
Xfanout509 net511 VSS VSS VCC VCC net509 sky130_fd_sc_hd__clkbuf_4
X_4292_ _1909_ _1919_ _1911_ _1910_ VSS VSS VCC VCC _1920_ sky130_fd_sc_hd__and4b_1
X_3243_ _0693_ _1185_ _0705_ VSS VSS VCC VCC _1187_ sky130_fd_sc_hd__a21o_1
X_3174_ _1129_ _1130_ net446 VSS VSS VCC VCC _1131_ sky130_fd_sc_hd__a21o_1
X_2958_ _0924_ _0926_ VSS VSS VCC VCC _0927_ sky130_fd_sc_hd__nor2_4
X_2889_ _0855_ _0856_ _0860_ _0807_ VSS VSS VCC VCC _0861_ sky130_fd_sc_hd__o2bb2a_1
X_4628_ net471 _2185_ _2186_ VSS VSS VCC VCC _2187_ sky130_fd_sc_hd__nor3_1
X_4559_ _2122_ _2114_ net716 VSS VSS VCC VCC _2124_ sky130_fd_sc_hd__o21ai_1
Xinput150 i_reg_data2[15] VSS VSS VCC VCC net150 sky130_fd_sc_hd__clkbuf_1
Xinput161 i_reg_data2[25] VSS VSS VCC VCC net161 sky130_fd_sc_hd__buf_2
Xinput172 i_reg_data2[6] VSS VSS VCC VCC net172 sky130_fd_sc_hd__clkbuf_1
X_3930_ net514 net244 net727 _1716_ VSS VSS VCC VCC _0093_ sky130_fd_sc_hd__o211a_1
X_3861_ net513 net87 net721 VSS VSS VCC VCC _1678_ sky130_fd_sc_hd__a21o_1
X_2812_ net671 u_bits.i_op2\[22\] _0784_ net349 VSS VSS VCC VCC _0786_ sky130_fd_sc_hd__o211a_1
X_3792_ net503 _1625_ VSS VSS VCC VCC _1626_ sky130_fd_sc_hd__and2b_1
X_2743_ net541 _0427_ _0457_ _0716_ VSS VSS VCC VCC _0718_ sky130_fd_sc_hd__o211ai_4
X_2674_ _0646_ _0648_ VSS VSS VCC VCC _0649_ sky130_fd_sc_hd__nand2_2
X_4413_ u_muldiv.o_div\[11\] _2028_ net471 net492 VSS VSS VCC VCC _2031_ sky130_fd_sc_hd__o2bb2a_1
X_4344_ _1970_ _1971_ _1969_ VSS VSS VCC VCC _1972_ sky130_fd_sc_hd__o21a_1
Xfanout317 _1993_ VSS VSS VCC VCC net317 sky130_fd_sc_hd__buf_6
Xfanout328 _0769_ VSS VSS VCC VCC net328 sky130_fd_sc_hd__buf_2
Xfanout339 net340 VSS VSS VCC VCC net339 sky130_fd_sc_hd__buf_4
X_4275_ u_muldiv.divisor\[15\] u_muldiv.dividend\[15\] VSS VSS VCC VCC _1903_
+ sky130_fd_sc_hd__and2b_1
X_3226_ _0614_ _0615_ _0625_ _1171_ VSS VSS VCC VCC _1174_ sky130_fd_sc_hd__a211o_1
X_3157_ _0810_ _0812_ _0982_ _1114_ net453 net450 VSS VSS VCC VCC _1115_ sky130_fd_sc_hd__mux4_2
X_3088_ net656 net658 net660 net662 net637 net625 VSS VSS VCC VCC _1050_ sky130_fd_sc_hd__mux4_1
X_4060_ net592 u_bits.i_op2\[14\] VSS VSS VCC VCC _1774_ sky130_fd_sc_hd__or2_1
X_3011_ net602 _0975_ net327 VSS VSS VCC VCC _0977_ sky130_fd_sc_hd__o21a_1
X_4962_ _1000_ _1001_ net407 VSS VSS VCC VCC _0406_ sky130_fd_sc_hd__and3_2
X_3913_ u_pc_sel.i_pc_next\[4\] net118 net390 VSS VSS VCC VCC _0079_ sky130_fd_sc_hd__mux2_1
X_4893_ u_muldiv.divisor\[0\] net498 net343 u_muldiv.divisor\[1\] vssd1 vssd1 vccd1
+ vccd1 _0345_ sky130_fd_sc_hd__a22o_1
X_3844_ net512 _1664_ VSS VSS VCC VCC _1665_ sky130_fd_sc_hd__and2b_1
X_3775_ net507 net237 net725 _1615_ VSS VSS VCC VCC _0039_ sky130_fd_sc_hd__o211a_1
X_2726_ net696 u_muldiv.add_prev\[11\] net542 VSS VSS VCC VCC _0701_ sky130_fd_sc_hd__mux2_1
X_2657_ _0614_ _0615_ VSS VSS VCC VCC _0632_ sky130_fd_sc_hd__nand2_1
X_5376_ clknet_leaf_159_i_clk _0403_ VSS VSS VCC VCC u_muldiv.mul\[55\] sky130_fd_sc_hd__dfxtp_1
X_2588_ net646 net555 net718 net537 net425 VSS VSS VCC VCC _0563_ sky130_fd_sc_hd__o2111ai_1
X_4327_ _1946_ _1947_ _1954_ VSS VSS VCC VCC _1955_ sky130_fd_sc_hd__and3_1
X_4258_ _0446_ u_muldiv.divisor\[10\] VSS VSS VCC VCC _1886_ sky130_fd_sc_hd__and2_1
X_3209_ u_pc_sel.i_inst_branch u_pc_sel.i_inst_jal_jalr VSS VSS VCC VCC net218
+ sky130_fd_sc_hd__or2_2
X_4189_ u_muldiv.mul\[19\] u_muldiv.mul\[18\] net404 VSS VSS VCC VCC _0233_
+ sky130_fd_sc_hd__mux2_1
Xfanout670 net671 VSS VSS VCC VCC net670 sky130_fd_sc_hd__buf_4
Xfanout681 u_bits.i_op1\[18\] VSS VSS VCC VCC net681 sky130_fd_sc_hd__buf_8
Xfanout692 u_bits.i_op1\[13\] VSS VSS VCC VCC net692 sky130_fd_sc_hd__buf_6
X_3560_ net528 _1445_ _1447_ _1448_ VSS VSS VCC VCC _1449_ sky130_fd_sc_hd__a2bb2o_1
X_2511_ net531 u_muldiv.add_prev\[20\] VSS VSS VCC VCC _0486_ sky130_fd_sc_hd__and2_1
X_3491_ _0425_ net569 net709 VSS VSS VCC VCC _1384_ sky130_fd_sc_hd__or3b_1
X_5230_ clknet_leaf_118_i_clk _0258_ VSS VSS VCC VCC u_muldiv.o_div\[7\] sky130_fd_sc_hd__dfxtp_2
X_2442_ u_muldiv.divisor\[2\] VSS VSS VCC VCC _0417_ sky130_fd_sc_hd__inv_2
X_5161_ clknet_leaf_76_i_clk _0193_ VSS VSS VCC VCC u_muldiv.add_prev\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_4112_ u_muldiv.divisor\[56\] net482 net337 u_muldiv.divisor\[57\] _1815_ vssd1 vssd1
+ vccd1 vccd1 _0176_ sky130_fd_sc_hd__a221o_1
X_5092_ clknet_leaf_50_i_clk _0125_ VSS VSS VCC VCC net308 sky130_fd_sc_hd__dfxtp_4
X_4043_ _1760_ net381 net594 VSS VSS VCC VCC _1761_ sky130_fd_sc_hd__a21oi_1
X_4945_ _1185_ _1189_ net406 VSS VSS VCC VCC _0389_ sky130_fd_sc_hd__and3_1
X_4876_ u_muldiv.dividend\[29\] u_muldiv.dividend\[28\] _2384_ u_muldiv.dividend\[30\]
+ VSS VSS VCC VCC _2413_ sky130_fd_sc_hd__o31a_1
X_3827_ net593 net595 net545 VSS VSS VCC VCC _1652_ sky130_fd_sc_hd__mux2_1
X_3758_ net666 net61 net389 VSS VSS VCC VCC _0027_ sky130_fd_sc_hd__mux2_1
X_2709_ _0669_ _0670_ _0680_ _0682_ VSS VSS VCC VCC _0684_ sky130_fd_sc_hd__nand4_4
X_3689_ net577 _1568_ VSS VSS VCC VCC _1569_ sky130_fd_sc_hd__nor2_1
Xoutput240 net504 VSS VSS VCC VCC o_ready sky130_fd_sc_hd__buf_2
Xoutput251 net251 VSS VSS VCC VCC o_result[15] sky130_fd_sc_hd__buf_2
Xoutput262 net262 VSS VSS VCC VCC o_result[25] sky130_fd_sc_hd__buf_2
Xoutput273 net273 VSS VSS VCC VCC o_result[6] sky130_fd_sc_hd__buf_2
X_5359_ clknet_leaf_85_i_clk _0386_ VSS VSS VCC VCC u_muldiv.mul\[38\] sky130_fd_sc_hd__dfxtp_2
Xoutput284 net284 VSS VSS VCC VCC o_wdata[14] sky130_fd_sc_hd__buf_2
Xoutput295 net295 VSS VSS VCC VCC o_wdata[24] sky130_fd_sc_hd__buf_2
X_2991_ net446 u_bits.i_op2\[26\] VSS VSS VCC VCC _0958_ sky130_fd_sc_hd__and2_1
X_4730_ u_muldiv.dividend\[15\] net462 u_muldiv.dividend\[16\] _2242_ vssd1 vssd1
+ vccd1 vccd1 _2280_ sky130_fd_sc_hd__nor4b_4
X_4661_ net695 _2215_ _2216_ VSS VSS VCC VCC _2217_ sky130_fd_sc_hd__o21ai_1
X_3612_ net573 net422 net345 _1082_ _1493_ VSS VSS VCC VCC _1497_ sky130_fd_sc_hd__a221o_1
X_4592_ _1865_ _1849_ _1850_ net459 VSS VSS VCC VCC _2154_ sky130_fd_sc_hd__a31o_1
X_3543_ net566 net556 u_muldiv.dividend\[8\] u_muldiv.mul\[40\] net362 vssd1 vssd1
+ vccd1 vccd1 _1433_ sky130_fd_sc_hd__a32o_1
X_3474_ net607 net614 net409 _1044_ VSS VSS VCC VCC _1368_ sky130_fd_sc_hd__or4_1
X_5213_ clknet_leaf_17_i_clk _0245_ VSS VSS VCC VCC u_muldiv.mul\[30\] sky130_fd_sc_hd__dfxtp_1
X_5144_ clknet_leaf_32_i_clk _0176_ VSS VSS VCC VCC u_muldiv.divisor\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_5075_ clknet_leaf_82_i_clk _0108_ VSS VSS VCC VCC net225 sky130_fd_sc_hd__dfxtp_4
X_4026_ net598 _1746_ _1747_ VSS VSS VCC VCC _1748_ sky130_fd_sc_hd__o21ba_1
X_4928_ u_muldiv.outsign net384 _2431_ _2430_ VSS VSS VCC VCC _0376_ sky130_fd_sc_hd__o22a_1
X_4859_ _2396_ _2397_ u_muldiv.dividend\[28\] net323 VSS VSS VCC VCC _0341_
+ sky130_fd_sc_hd__a2bb2o_1
X_3190_ net651 u_bits.i_op2\[31\] VSS VSS VCC VCC _1146_ sky130_fd_sc_hd__nand2_1
X_2974_ net690 net693 net695 net697 net642 net630 VSS VSS VCC VCC _0942_ sky130_fd_sc_hd__mux4_2
X_4713_ _1908_ _1915_ _0413_ VSS VSS VCC VCC _2264_ sky130_fd_sc_hd__a21oi_1
X_4644_ u_muldiv.dividend\[10\] u_muldiv.dividend\[9\] _2180_ VSS VSS VCC VCC
+ _2201_ sky130_fd_sc_hd__or3_2
X_4575_ net438 _2136_ _2138_ _2135_ VSS VSS VCC VCC _2139_ sky130_fd_sc_hd__o31ai_1
X_3526_ _0426_ _0436_ net573 net421 VSS VSS VCC VCC _1417_ sky130_fd_sc_hd__o211a_1
X_3457_ _0422_ _1350_ _1351_ net354 net208 VSS VSS VCC VCC _1352_ sky130_fd_sc_hd__a32o_1
X_3388_ net572 net421 _0846_ net520 VSS VSS VCC VCC _1286_ sky130_fd_sc_hd__a31o_1
X_5127_ clknet_4_4__leaf_i_clk _0159_ VSS VSS VCC VCC u_muldiv.divisor\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_5058_ clknet_leaf_30_i_clk _0091_ VSS VSS VCC VCC net242 sky130_fd_sc_hd__dfxtp_4
X_4009_ net640 net626 net346 net378 VSS VSS VCC VCC _1734_ sky130_fd_sc_hd__o31a_1
X_2690_ _0663_ _0664_ net428 VSS VSS VCC VCC _0665_ sky130_fd_sc_hd__a21o_1
X_4360_ _1987_ VSS VSS VCC VCC _1988_ sky130_fd_sc_hd__clkinv_2
X_3311_ _1128_ _1132_ u_adder.i_cmp_inverse VSS VSS VCC VCC _1241_ sky130_fd_sc_hd__a21oi_1
X_4291_ _1915_ _1916_ _1918_ VSS VSS VCC VCC _1919_ sky130_fd_sc_hd__and3_1
X_3242_ _0693_ _0705_ _1185_ VSS VSS VCC VCC _1186_ sky130_fd_sc_hd__nand3_2
X_3173_ _0459_ net423 net651 _0781_ VSS VSS VCC VCC _1130_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_121_i_clk clknet_4_11__leaf_i_clk VSS VSS VCC VCC clknet_leaf_121_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2957_ _0922_ _0923_ VSS VSS VCC VCC _0926_ sky130_fd_sc_hd__nor2_1
X_2888_ _0858_ _0859_ net623 VSS VSS VCC VCC _0860_ sky130_fd_sc_hd__mux2_1
X_4627_ _2184_ net373 net702 VSS VSS VCC VCC _2186_ sky130_fd_sc_hd__and3_1
X_4558_ net716 _2122_ _2114_ VSS VSS VCC VCC _2123_ sky130_fd_sc_hd__or3_1
X_3509_ u_bits.i_op2\[6\] net706 _1400_ net350 VSS VSS VCC VCC _1401_ sky130_fd_sc_hd__o211ai_1
X_4489_ u_muldiv.o_div\[27\] _2088_ net475 net465 VSS VSS VCC VCC _2091_ sky130_fd_sc_hd__o2bb2a_1
Xinput140 i_rd[1] VSS VSS VCC VCC net140 sky130_fd_sc_hd__clkbuf_2
Xinput151 i_reg_data2[16] VSS VSS VCC VCC net151 sky130_fd_sc_hd__clkbuf_1
Xinput162 i_reg_data2[26] VSS VSS VCC VCC net162 sky130_fd_sc_hd__clkbuf_1
Xinput173 i_reg_data2[7] VSS VSS VCC VCC net173 sky130_fd_sc_hd__clkbuf_1
X_3860_ net512 _1676_ VSS VSS VCC VCC _1677_ sky130_fd_sc_hd__and2b_1
X_2811_ net570 net440 VSS VSS VCC VCC _0785_ sky130_fd_sc_hd__nor2_4
X_3791_ net618 net626 net545 VSS VSS VCC VCC _1625_ sky130_fd_sc_hd__mux2_1
X_2742_ net541 _0427_ _0716_ VSS VSS VCC VCC _0717_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_4_11__f_i_clk clknet_2_2_0_i_clk VSS VSS VCC VCC clknet_4_11__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_2673_ _0644_ _0647_ VSS VSS VCC VCC _0648_ sky130_fd_sc_hd__nand2_2
X_4412_ u_muldiv.o_div\[10\] net331 net375 net318 _2030_ VSS VSS VCC VCC _0261_
+ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_68_i_clk clknet_4_13__leaf_i_clk VSS VSS VCC VCC clknet_leaf_68_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_4343_ u_muldiv.divisor\[30\] u_muldiv.dividend\[30\] VSS VSS VCC VCC _1971_
+ sky130_fd_sc_hd__and2_1
Xfanout318 net319 VSS VSS VCC VCC net318 sky130_fd_sc_hd__buf_4
Xfanout329 net330 VSS VSS VCC VCC net329 sky130_fd_sc_hd__clkbuf_8
X_4274_ u_muldiv.divisor\[14\] u_muldiv.dividend\[14\] VSS VSS VCC VCC _1902_
+ sky130_fd_sc_hd__xor2_1
X_3225_ _0625_ _1171_ _0614_ _0615_ VSS VSS VCC VCC _1173_ sky130_fd_sc_hd__o211ai_4
X_3156_ net652 net654 net656 net658 net638 net627 VSS VSS VCC VCC _1114_ sky130_fd_sc_hd__mux4_1
X_3087_ net620 _0902_ _1048_ VSS VSS VCC VCC _1049_ sky130_fd_sc_hd__a21o_2
X_3989_ net43 net40 net391 _1718_ VSS VSS VCC VCC _0150_ sky130_fd_sc_hd__a31o_1
X_3010_ net612 _0974_ net347 VSS VSS VCC VCC _0976_ sky130_fd_sc_hd__o21ai_1
X_4961_ _0970_ net400 VSS VSS VCC VCC _0405_ sky130_fd_sc_hd__nor2_2
X_3912_ u_pc_sel.i_pc_next\[3\] net117 net398 VSS VSS VCC VCC _0078_ sky130_fd_sc_hd__mux2_1
X_4892_ u_muldiv.dividend\[31\] net323 _2424_ _2427_ VSS VSS VCC VCC _0344_
+ sky130_fd_sc_hd__o2bb2ai_1
X_3843_ net590 u_bits.i_op2\[14\] net548 VSS VSS VCC VCC _1664_ sky130_fd_sc_hd__mux2_1
X_3774_ net141 net507 VSS VSS VCC VCC _1615_ sky130_fd_sc_hd__nand2b_1
X_2725_ _0696_ _0697_ net429 VSS VSS VCC VCC _0700_ sky130_fd_sc_hd__a21oi_2
X_2656_ _0620_ _0621_ _0624_ VSS VSS VCC VCC _0631_ sky130_fd_sc_hd__nand3_1
X_2587_ _0554_ _0561_ _0560_ VSS VSS VCC VCC _0562_ sky130_fd_sc_hd__o21a_1
X_5375_ clknet_leaf_159_i_clk _0402_ VSS VSS VCC VCC u_muldiv.mul\[54\] sky130_fd_sc_hd__dfxtp_1
X_4326_ _1948_ _1949_ _1951_ _1952_ VSS VSS VCC VCC _1954_ sky130_fd_sc_hd__and4_1
X_4257_ u_muldiv.divisor\[10\] _0446_ VSS VSS VCC VCC _1885_ sky130_fd_sc_hd__nor2_1
X_3208_ net514 net563 _1161_ net499 VSS VSS VCC VCC mul_op2_signed_next sky130_fd_sc_hd__and4bb_1
X_4188_ u_muldiv.mul\[18\] u_muldiv.mul\[17\] net404 VSS VSS VCC VCC _0232_
+ sky130_fd_sc_hd__mux2_1
X_3139_ _1097_ VSS VSS VCC VCC _1098_ sky130_fd_sc_hd__inv_2
Xfanout660 u_bits.i_op1\[26\] VSS VSS VCC VCC net660 sky130_fd_sc_hd__buf_4
Xfanout671 u_bits.i_op1\[22\] VSS VSS VCC VCC net671 sky130_fd_sc_hd__buf_8
Xfanout682 net683 VSS VSS VCC VCC net682 sky130_fd_sc_hd__buf_6
Xfanout693 net694 VSS VSS VCC VCC net693 sky130_fd_sc_hd__buf_6
X_2510_ _0483_ net432 VSS VSS VCC VCC _0485_ sky130_fd_sc_hd__nand2_1
X_3490_ net609 net617 net409 _1081_ VSS VSS VCC VCC _1383_ sky130_fd_sc_hd__or4_1
X_2441_ u_muldiv.divisor\[11\] VSS VSS VCC VCC _0416_ sky130_fd_sc_hd__inv_2
X_5160_ clknet_leaf_75_i_clk _0192_ VSS VSS VCC VCC u_muldiv.add_prev\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_4111_ net584 _1813_ _1814_ VSS VSS VCC VCC _1815_ sky130_fd_sc_hd__a21oi_1
X_5091_ clknet_leaf_164_i_clk _0124_ VSS VSS VCC VCC net307 sky130_fd_sc_hd__dfxtp_4
X_4042_ net597 net596 net595 _1749_ VSS VSS VCC VCC _1760_ sky130_fd_sc_hd__or4_2
X_4944_ _1179_ _1180_ net406 VSS VSS VCC VCC _0388_ sky130_fd_sc_hd__and3_1
X_4875_ u_muldiv.dividend\[30\] _2402_ VSS VSS VCC VCC _2412_ sky130_fd_sc_hd__nor2_1
X_3826_ net595 net724 _1651_ _1650_ VSS VSS VCC VCC _0054_ sky130_fd_sc_hd__o22a_1
X_3757_ net669 net60 net392 VSS VSS VCC VCC _0026_ sky130_fd_sc_hd__mux2_1
X_2708_ _0680_ _0682_ VSS VSS VCC VCC _0683_ sky130_fd_sc_hd__nand2_1
X_3688_ _1558_ _1567_ net733 VSS VSS VCC VCC _1568_ sky130_fd_sc_hd__a21oi_4
Xoutput230 net230 VSS VSS VCC VCC o_pc_target[5] sky130_fd_sc_hd__buf_2
X_2639_ _0609_ _0610_ _0613_ VSS VSS VCC VCC _0614_ sky130_fd_sc_hd__nand3_2
Xoutput241 net241 VSS VSS VCC VCC o_reg_write sky130_fd_sc_hd__buf_2
Xoutput252 net252 VSS VSS VCC VCC o_result[16] sky130_fd_sc_hd__buf_2
Xoutput263 net263 VSS VSS VCC VCC o_result[26] sky130_fd_sc_hd__buf_2
Xoutput274 net274 VSS VSS VCC VCC o_result[7] sky130_fd_sc_hd__buf_2
X_5358_ clknet_leaf_86_i_clk _0385_ VSS VSS VCC VCC u_muldiv.mul\[37\] sky130_fd_sc_hd__dfxtp_1
Xoutput285 net285 VSS VSS VCC VCC o_wdata[15] sky130_fd_sc_hd__buf_2
Xoutput296 net296 VSS VSS VCC VCC o_wdata[25] sky130_fd_sc_hd__buf_2
X_4309_ u_muldiv.dividend\[21\] u_muldiv.divisor\[21\] VSS VSS VCC VCC _1937_
+ sky130_fd_sc_hd__and2b_1
X_5289_ clknet_4_14__leaf_i_clk _0317_ VSS VSS VCC VCC u_muldiv.dividend\[4\]
+ sky130_fd_sc_hd__dfxtp_2
Xfanout490 net495 VSS VSS VCC VCC net490 sky130_fd_sc_hd__buf_4
X_2990_ net729 _0956_ _0957_ net574 VSS VSS VCC VCC net262 sky130_fd_sc_hd__a211oi_4
X_4660_ _2215_ net695 net472 VSS VSS VCC VCC _2216_ sky130_fd_sc_hd__a21oi_1
X_3611_ net604 _1495_ net364 net573 VSS VSS VCC VCC _1496_ sky130_fd_sc_hd__o211a_1
X_4591_ _1850_ _1865_ _1849_ VSS VSS VCC VCC _2153_ sky130_fd_sc_hd__a21oi_1
X_3542_ net520 _1431_ net354 net213 VSS VSS VCC VCC _1432_ sky130_fd_sc_hd__a2bb2o_1
X_3473_ net604 _1361_ _1366_ net573 net365 VSS VSS VCC VCC _1367_ sky130_fd_sc_hd__o2111ai_4
X_5212_ clknet_leaf_19_i_clk _0244_ VSS VSS VCC VCC u_muldiv.mul\[29\] sky130_fd_sc_hd__dfxtp_1
X_5143_ clknet_leaf_32_i_clk _0175_ VSS VSS VCC VCC u_muldiv.divisor\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_5074_ clknet_leaf_81_i_clk _0107_ VSS VSS VCC VCC net224 sky130_fd_sc_hd__dfxtp_1
X_4025_ _1745_ net379 net598 net329 VSS VSS VCC VCC _1747_ sky130_fd_sc_hd__a31o_1
X_4927_ net651 _1266_ net487 net468 VSS VSS VCC VCC _2431_ sky130_fd_sc_hd__a211o_1
X_4858_ net476 _2393_ net315 VSS VSS VCC VCC _2397_ sky130_fd_sc_hd__o21ai_1
X_3809_ net505 net105 net719 VSS VSS VCC VCC _1639_ sky130_fd_sc_hd__a21o_1
X_4789_ _2333_ _2325_ net480 _2332_ VSS VSS VCC VCC _2334_ sky130_fd_sc_hd__o22ai_1
X_2973_ net628 _0897_ _0847_ net613 _0940_ VSS VSS VCC VCC _0941_ sky130_fd_sc_hd__o32a_1
X_4712_ _2261_ _2262_ net437 VSS VSS VCC VCC _2263_ sky130_fd_sc_hd__a21o_1
X_4643_ u_muldiv.dividend\[9\] _2180_ u_muldiv.dividend\[10\] VSS VSS VCC VCC
+ _2200_ sky130_fd_sc_hd__o21ai_1
X_4574_ u_muldiv.dividend\[0\] net464 u_muldiv.dividend\[2\] u_muldiv.dividend\[3\]
+ VSS VSS VCC VCC _2138_ sky130_fd_sc_hd__o31a_1
X_3525_ _1412_ _0765_ _1415_ VSS VSS VCC VCC _1416_ sky130_fd_sc_hd__a21boi_2
X_3456_ net617 net712 _0781_ net441 VSS VSS VCC VCC _1351_ sky130_fd_sc_hd__a211o_1
X_3387_ _0765_ _1278_ _1284_ VSS VSS VCC VCC _1285_ sky130_fd_sc_hd__a21oi_2
X_5126_ clknet_leaf_28_i_clk _0158_ VSS VSS VCC VCC u_muldiv.divisor\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_5057_ clknet_leaf_47_i_clk _0090_ VSS VSS VCC VCC u_pc_sel.i_pc_next\[15\]
+ sky130_fd_sc_hd__dfxtp_4
X_4008_ u_muldiv.divisor\[34\] net478 net333 u_muldiv.divisor\[35\] _1733_ vssd1 vssd1
+ vccd1 vccd1 _0154_ sky130_fd_sc_hd__a221o_1
Xclkbuf_4_9__f_i_clk clknet_2_2_0_i_clk VSS VSS VCC VCC clknet_4_9__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_3310_ _1238_ _1239_ u_adder.i_cmp_inverse VSS VSS VCC VCC _1240_ sky130_fd_sc_hd__a21boi_1
X_4290_ net462 u_muldiv.divisor\[17\] VSS VSS VCC VCC _1918_ sky130_fd_sc_hd__nand2b_1
X_3241_ _0733_ _1184_ _0695_ VSS VSS VCC VCC _1185_ sky130_fd_sc_hd__o21ai_4
X_3172_ net641 net549 net651 _0781_ net423 VSS VSS VCC VCC _1129_ sky130_fd_sc_hd__o2111ai_1
X_2956_ _0922_ _0923_ VSS VSS VCC VCC _0925_ sky130_fd_sc_hd__nand2_1
X_2887_ net678 net681 u_bits.i_op1\[17\] net685 net639 net634 VSS VSS VCC VCC
+ _0859_ sky130_fd_sc_hd__mux4_1
X_4626_ _2184_ net373 net702 VSS VSS VCC VCC _2185_ sky130_fd_sc_hd__a21oi_1
X_4557_ net461 net718 VSS VSS VCC VCC _2122_ sky130_fd_sc_hd__nor2_1
X_3508_ net568 net706 u_bits.i_op2\[6\] VSS VSS VCC VCC _1400_ sky130_fd_sc_hd__nand3b_1
X_4488_ u_muldiv.o_div\[26\] net330 _1991_ net315 _2090_ VSS VSS VCC VCC _0277_
+ sky130_fd_sc_hd__a32o_1
X_3439_ net443 _1331_ _1334_ net733 VSS VSS VCC VCC _1335_ sky130_fd_sc_hd__a211o_2
X_5109_ clknet_leaf_43_i_clk _0142_ VSS VSS VCC VCC u_wr_mux.i_reg_data2\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput130 i_pc_target[1] VSS VSS VCC VCC net130 sky130_fd_sc_hd__clkbuf_8
Xinput141 i_rd[2] VSS VSS VCC VCC net141 sky130_fd_sc_hd__buf_6
Xinput152 i_reg_data2[17] VSS VSS VCC VCC net152 sky130_fd_sc_hd__clkbuf_1
Xinput163 i_reg_data2[27] VSS VSS VCC VCC net163 sky130_fd_sc_hd__clkbuf_1
Xinput174 i_reg_data2[8] VSS VSS VCC VCC net174 sky130_fd_sc_hd__clkbuf_1
X_2810_ net564 u_bits.i_op2\[22\] u_bits.i_op1\[22\] VSS VSS VCC VCC _0784_
+ sky130_fd_sc_hd__nand3b_1
X_3790_ net636 net727 _1624_ _1623_ VSS VSS VCC VCC _0045_ sky130_fd_sc_hd__o22a_1
X_2741_ net648 net554 net700 net541 net425 VSS VSS VCC VCC _0716_ sky130_fd_sc_hd__o2111ai_4
X_2672_ net428 _0640_ _0641_ _0645_ VSS VSS VCC VCC _0647_ sky130_fd_sc_hd__a31oi_1
X_4411_ net470 u_muldiv.quotient_msk\[10\] net435 _2028_ _2029_ vssd1 vssd1 vccd1
+ vccd1 _2030_ sky130_fd_sc_hd__a32o_1
X_4342_ u_muldiv.divisor\[30\] u_muldiv.dividend\[30\] VSS VSS VCC VCC _1970_
+ sky130_fd_sc_hd__nor2_2
Xfanout319 net321 VSS VSS VCC VCC net319 sky130_fd_sc_hd__clkbuf_8
X_4273_ _1893_ _1898_ _1900_ VSS VSS VCC VCC _1901_ sky130_fd_sc_hd__a21oi_2
X_3224_ _0606_ _0629_ _0633_ VSS VSS VCC VCC _1172_ sky130_fd_sc_hd__a21o_1
