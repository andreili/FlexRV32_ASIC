* NGSPICE file created from rv_decode.ext - technology: sky130A

.ends

.ends

.ends

.ends

.ends

.ends

.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt rv_decode i_clk i_flush i_instruction[0] i_instruction[10] i_instruction[11]
+ i_instruction[12] i_instruction[13] i_instruction[14] i_instruction[15] i_instruction[16]
+ i_instruction[17] i_instruction[18] i_instruction[19] i_instruction[1] i_instruction[20]
+ i_instruction[21] i_instruction[22] i_instruction[23] i_instruction[24] i_instruction[25]
+ i_instruction[26] i_instruction[27] i_instruction[28] i_instruction[29] i_instruction[2]
+ i_instruction[30] i_instruction[31] i_instruction[3] i_instruction[4] i_instruction[5]
+ i_instruction[6] i_instruction[7] i_instruction[8] i_instruction[9] i_pc[10] i_pc[11]
+ i_pc[12] i_pc[13] i_pc[14] i_pc[15] i_pc[1] i_pc[2] i_pc[3] i_pc[4] i_pc[5] i_pc[6]
+ i_pc[7] i_pc[8] i_pc[9] i_pc_next[10] i_pc_next[11] i_pc_next[12] i_pc_next[13]
+ i_pc_next[14] i_pc_next[15] i_pc_next[1] i_pc_next[2] i_pc_next[3] i_pc_next[4]
+ i_pc_next[5] i_pc_next[6] i_pc_next[7] i_pc_next[8] i_pc_next[9] i_ready i_stall
+ o_alu_ctrl[0] o_alu_ctrl[1] o_alu_ctrl[2] o_alu_ctrl[3] o_alu_ctrl[4] o_csr_clear
+ o_csr_ebreak o_csr_idx[0] o_csr_idx[10] o_csr_idx[11] o_csr_idx[1] o_csr_idx[2]
+ o_csr_idx[3] o_csr_idx[4] o_csr_idx[5] o_csr_idx[6] o_csr_idx[7] o_csr_idx[8] o_csr_idx[9]
+ o_csr_imm[0] o_csr_imm[1] o_csr_imm[2] o_csr_imm[3] o_csr_imm[4] o_csr_imm_sel o_csr_read
+ o_csr_set o_csr_write o_funct3[0] o_funct3[1] o_funct3[2] o_imm_i[0] o_imm_i[10]
+ o_imm_i[11] o_imm_i[12] o_imm_i[13] o_imm_i[14] o_imm_i[15] o_imm_i[16] o_imm_i[17]
+ o_imm_i[18] o_imm_i[19] o_imm_i[1] o_imm_i[20] o_imm_i[21] o_imm_i[22] o_imm_i[23]
+ o_imm_i[24] o_imm_i[25] o_imm_i[26] o_imm_i[27] o_imm_i[28] o_imm_i[29] o_imm_i[2]
+ o_imm_i[30] o_imm_i[31] o_imm_i[3] o_imm_i[4] o_imm_i[5] o_imm_i[6] o_imm_i[7] o_imm_i[8]
+ o_imm_i[9] o_inst_branch o_inst_jal o_inst_jalr o_inst_mret o_inst_store o_inst_supported
+ o_op1_src o_op2_src o_pc[10] o_pc[11] o_pc[12] o_pc[13] o_pc[14] o_pc[15] o_pc[1]
+ o_pc[2] o_pc[3] o_pc[4] o_pc[5] o_pc[6] o_pc[7] o_pc[8] o_pc[9] o_pc_next[10] o_pc_next[11]
+ o_pc_next[12] o_pc_next[13] o_pc_next[14] o_pc_next[15] o_pc_next[1] o_pc_next[2]
+ o_pc_next[3] o_pc_next[4] o_pc_next[5] o_pc_next[6] o_pc_next[7] o_pc_next[8] o_pc_next[9]
+ o_rd[0] o_rd[1] o_rd[2] o_rd[3] o_rd[4] o_reg_write o_res_src[0] o_res_src[1] o_res_src[2]
+ o_rs1[0] o_rs1[1] o_rs1[2] o_rs1[3] o_rs1[4] o_rs2[0] o_rs2[1] o_rs2[2] o_rs2[3]
+ o_rs2[4] vccd1 vssd1
X_501_ o_pc_next[6] i_pc_next[6] net21 vssd1 vssd1 vccd1 vccd1 _005_ sky130_fd_sc_hd__mux2_1
X_432_ o_rd[0] o_inst_store _092_ o_csr_idx[0] vssd1 vssd1 vccd1 vccd1 _093_ sky130_fd_sc_hd__a22o_1
X_415_ o_res_src[1] o_res_src[2] vssd1 vssd1 vccd1 vccd1 o_res_src[0] sky130_fd_sc_hd__nor2_4
X_895_ o_csr_imm_sel vssd1 vssd1 vccd1 vccd1 o_funct3[2] sky130_fd_sc_hd__buf_2
X_680_ net28 o_csr_imm[0] net25 _267_ vssd1 vssd1 vccd1 vccd1 _031_ sky130_fd_sc_hd__o211a_2
X_878_ clknet_3_7__leaf_i_clk _047_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[11] sky130_fd_sc_hd__dfxtp_4
Xfanout7 _159_ vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_4
X_801_ _373_ _374_ _375_ net12 net30 vssd1 vssd1 vccd1 vccd1 _376_ sky130_fd_sc_hd__a221o_1
X_732_ net28 o_csr_idx[1] _311_ _313_ net25 vssd1 vssd1 vccd1 vccd1 _037_ sky130_fd_sc_hd__o221a_4
X_663_ net26 o_funct3[1] _249_ _252_ net23 vssd1 vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__o221a_1
X_594_ net43 _165_ vssd1 vssd1 vccd1 vccd1 _192_ sky130_fd_sc_hd__or2_1
X_715_ _128_ _130_ _154_ vssd1 vssd1 vccd1 vccd1 _298_ sky130_fd_sc_hd__or3b_1
X_646_ net26 o_rd[4] net23 _237_ vssd1 vssd1 vccd1 vccd1 _027_ sky130_fd_sc_hd__o211a_1
X_577_ i_instruction[3] _173_ _171_ vssd1 vssd1 vccd1 vccd1 _177_ sky130_fd_sc_hd__a21bo_1
X_500_ o_pc_next[5] i_pc_next[5] net22 vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__mux2_2
X_431_ _090_ _091_ vssd1 vssd1 vccd1 vccd1 _092_ sky130_fd_sc_hd__and2_4
X_629_ net27 o_rd[1] vssd1 vssd1 vccd1 vccd1 _224_ sky130_fd_sc_hd__or2_1
X_414_ instruction\[5\] instruction\[1\] instruction\[0\] _083_ vssd1 vssd1 vccd1
+ vccd1 o_res_src[2] sky130_fd_sc_hd__and4b_4
X_894_ o_alu_ctrl[3] vssd1 vssd1 vccd1 vccd1 o_csr_idx[10] sky130_fd_sc_hd__buf_2
X_877_ clknet_3_4__leaf_i_clk _046_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[3] sky130_fd_sc_hd__dfxtp_4
Xfanout8 _144_ vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_4
X_800_ net34 i_instruction[9] _120_ net8 i_instruction[28] vssd1 vssd1 vccd1 vccd1
+ _375_ sky130_fd_sc_hd__a32o_1
X_731_ net18 net12 _312_ net30 vssd1 vssd1 vccd1 vccd1 _313_ sky130_fd_sc_hd__a31o_1
X_662_ _188_ _250_ _251_ net29 vssd1 vssd1 vccd1 vccd1 _252_ sky130_fd_sc_hd__a211o_1
X_593_ _166_ _190_ _189_ _168_ vssd1 vssd1 vccd1 vccd1 _191_ sky130_fd_sc_hd__o211ai_1
X_714_ net8 _150_ vssd1 vssd1 vccd1 vccd1 _297_ sky130_fd_sc_hd__nor2_1
X_645_ _123_ _158_ _235_ _236_ net30 vssd1 vssd1 vccd1 vccd1 _237_ sky130_fd_sc_hd__a41o_1
X_576_ i_flush _176_ vssd1 vssd1 vccd1 vccd1 _018_ sky130_fd_sc_hd__nor2_1
X_430_ instruction\[3\] _084_ instruction\[2\] _077_ vssd1 vssd1 vccd1 vccd1 _091_
+ sky130_fd_sc_hd__or4b_2
X_628_ _216_ _217_ _222_ net13 vssd1 vssd1 vccd1 vccd1 _223_ sky130_fd_sc_hd__o22a_1
X_559_ i_instruction[1] _136_ vssd1 vssd1 vccd1 vccd1 _160_ sky130_fd_sc_hd__or2_4
X_413_ instruction\[1\] instruction\[0\] vssd1 vssd1 vccd1 vccd1 _084_ sky130_fd_sc_hd__nand2_4
X_893_ clknet_3_3__leaf_i_clk _062_ vssd1 vssd1 vccd1 vccd1 o_pc[15] sky130_fd_sc_hd__dfxtp_2
X_876_ clknet_3_4__leaf_i_clk _045_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[9] sky130_fd_sc_hd__dfxtp_4
Xfanout9 _144_ vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_2
X_730_ i_instruction[21] _152_ _145_ vssd1 vssd1 vccd1 vccd1 _312_ sky130_fd_sc_hd__mux2_1
X_661_ net43 _135_ _137_ _183_ vssd1 vssd1 vccd1 vccd1 _251_ sky130_fd_sc_hd__a31o_1
X_592_ i_instruction[10] _123_ vssd1 vssd1 vccd1 vccd1 _190_ sky130_fd_sc_hd__nand2_1
X_859_ clknet_3_5__leaf_i_clk _028_ vssd1 vssd1 vccd1 vccd1 o_funct3[0] sky130_fd_sc_hd__dfxtp_4
X_713_ i_flush _296_ vssd1 vssd1 vccd1 vccd1 _035_ sky130_fd_sc_hd__nor2_1
X_644_ _075_ net12 vssd1 vssd1 vccd1 vccd1 _236_ sky130_fd_sc_hd__nand2_1
X_575_ net31 instruction\[2\] _174_ _175_ vssd1 vssd1 vccd1 vccd1 _176_ sky130_fd_sc_hd__o2bb2a_1
X_627_ _157_ _221_ _220_ _138_ vssd1 vssd1 vccd1 vccd1 _222_ sky130_fd_sc_hd__a2bb2o_1
X_558_ i_instruction[1] _136_ vssd1 vssd1 vccd1 vccd1 _159_ sky130_fd_sc_hd__nor2_4
X_489_ _067_ instruction\[2\] instruction\[3\] instruction\[6\] vssd1 vssd1 vccd1
+ vccd1 _109_ sky130_fd_sc_hd__a211o_1
X_412_ _066_ _067_ _068_ vssd1 vssd1 vccd1 vccd1 _083_ sky130_fd_sc_hd__and3_2
X_892_ clknet_3_2__leaf_i_clk _061_ vssd1 vssd1 vccd1 vccd1 o_pc[14] sky130_fd_sc_hd__dfxtp_2
X_875_ clknet_3_4__leaf_i_clk _044_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[8] sky130_fd_sc_hd__dfxtp_4
X_660_ _120_ net10 vssd1 vssd1 vccd1 vccd1 _250_ sky130_fd_sc_hd__nor2_2
X_591_ _166_ _187_ vssd1 vssd1 vccd1 vccd1 _189_ sky130_fd_sc_hd__or2_1
X_858_ clknet_3_5__leaf_i_clk _027_ vssd1 vssd1 vccd1 vccd1 o_rd[4] sky130_fd_sc_hd__dfxtp_2
X_789_ _243_ _364_ i_instruction[27] _172_ vssd1 vssd1 vccd1 vccd1 _365_ sky130_fd_sc_hd__a2bb2o_1
X_712_ net29 o_csr_imm[4] _295_ vssd1 vssd1 vccd1 vccd1 _296_ sky130_fd_sc_hd__a21oi_1
X_643_ net19 net5 _193_ vssd1 vssd1 vccd1 vccd1 _235_ sky130_fd_sc_hd__or3_1
X_574_ net6 _168_ _170_ _146_ vssd1 vssd1 vccd1 vccd1 _175_ sky130_fd_sc_hd__a31o_1
X_626_ _145_ _156_ _159_ _127_ vssd1 vssd1 vccd1 vccd1 _221_ sky130_fd_sc_hd__a211o_1
X_557_ _118_ _157_ vssd1 vssd1 vccd1 vccd1 _158_ sky130_fd_sc_hd__nand2_4
X_488_ o_csr_imm_sel o_funct3[1] instruction\[6\] instruction\[5\] vssd1 vssd1 vccd1
+ vccd1 _108_ sky130_fd_sc_hd__or4_1
X_411_ o_inst_branch _081_ _082_ vssd1 vssd1 vccd1 vccd1 o_op2_src sky130_fd_sc_hd__nor3_4
X_609_ i_instruction[7] _129_ _204_ vssd1 vssd1 vccd1 vccd1 _205_ sky130_fd_sc_hd__mux2_1
X_891_ clknet_3_5__leaf_i_clk _060_ vssd1 vssd1 vccd1 vccd1 o_pc[13] sky130_fd_sc_hd__dfxtp_2
X_874_ clknet_3_6__leaf_i_clk _043_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[7] sky130_fd_sc_hd__dfxtp_4
X_590_ net43 _145_ vssd1 vssd1 vccd1 vccd1 _188_ sky130_fd_sc_hd__or2_4
X_857_ clknet_3_7__leaf_i_clk _026_ vssd1 vssd1 vccd1 vccd1 o_rd[3] sky130_fd_sc_hd__dfxtp_2
X_788_ i_instruction[3] _164_ _363_ vssd1 vssd1 vccd1 vccd1 _364_ sky130_fd_sc_hd__a21oi_1
X_711_ net5 _294_ _292_ _147_ vssd1 vssd1 vccd1 vccd1 _295_ sky130_fd_sc_hd__o211a_2
X_642_ net26 o_rd[3] net23 _233_ _234_ vssd1 vssd1 vccd1 vccd1 _026_ sky130_fd_sc_hd__o2111a_1
X_573_ _150_ net14 _158_ _161_ net5 vssd1 vssd1 vccd1 vccd1 _174_ sky130_fd_sc_hd__o221a_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_625_ _121_ _218_ _219_ _126_ _193_ vssd1 vssd1 vccd1 vccd1 _220_ sky130_fd_sc_hd__a32o_1
X_556_ _154_ _156_ vssd1 vssd1 vccd1 vccd1 _157_ sky130_fd_sc_hd__and2_1
X_487_ instruction\[5\] _067_ _076_ _084_ vssd1 vssd1 vccd1 vccd1 o_reg_write sky130_fd_sc_hd__a31oi_4
X_410_ instruction\[5\] instruction\[4\] _076_ instruction\[6\] vssd1 vssd1 vccd1
+ vccd1 _082_ sky130_fd_sc_hd__and4b_1
X_608_ _164_ _187_ vssd1 vssd1 vccd1 vccd1 _204_ sky130_fd_sc_hd__nor2_1
X_539_ _116_ _141_ i_flush vssd1 vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__a21oi_1
X_890_ clknet_3_2__leaf_i_clk _059_ vssd1 vssd1 vccd1 vccd1 o_pc[12] sky130_fd_sc_hd__dfxtp_2
X_873_ clknet_3_7__leaf_i_clk _042_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[6] sky130_fd_sc_hd__dfxtp_2
X_856_ clknet_3_3__leaf_i_clk _025_ vssd1 vssd1 vccd1 vccd1 o_rd[2] sky130_fd_sc_hd__dfxtp_2
X_787_ _126_ _145_ _165_ vssd1 vssd1 vccd1 vccd1 _363_ sky130_fd_sc_hd__and3_1
X_710_ _123_ _195_ _257_ _293_ vssd1 vssd1 vccd1 vccd1 _294_ sky130_fd_sc_hd__a211o_1
X_641_ net31 _122_ net10 _225_ vssd1 vssd1 vccd1 vccd1 _234_ sky130_fd_sc_hd__or4_1
X_572_ net5 _172_ vssd1 vssd1 vccd1 vccd1 _173_ sky130_fd_sc_hd__and2_4
X_839_ clknet_3_7__leaf_i_clk _008_ vssd1 vssd1 vccd1 vccd1 o_pc_next[9] sky130_fd_sc_hd__dfxtp_2
X_624_ _152_ i_instruction[8] _189_ vssd1 vssd1 vccd1 vccd1 _219_ sky130_fd_sc_hd__mux2_1
X_555_ net40 net14 vssd1 vssd1 vccd1 vccd1 _156_ sky130_fd_sc_hd__and2_1
X_486_ o_funct3[1] o_funct3[0] _085_ vssd1 vssd1 vccd1 vccd1 o_csr_clear sky130_fd_sc_hd__and3_2
X_607_ _201_ _203_ i_flush vssd1 vssd1 vccd1 vccd1 _022_ sky130_fd_sc_hd__a21oi_1
X_538_ _118_ _134_ net13 net31 vssd1 vssd1 vccd1 vccd1 _141_ sky130_fd_sc_hd__a31o_1
X_469_ o_csr_idx[7] net4 net1 vssd1 vssd1 vccd1 vccd1 o_imm_i[27] sky130_fd_sc_hd__a21o_2
Xclkbuf_3_2__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_872_ clknet_3_5__leaf_i_clk _041_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[5] sky130_fd_sc_hd__dfxtp_4
X_855_ clknet_3_0__leaf_i_clk _024_ vssd1 vssd1 vccd1 vccd1 o_rd[1] sky130_fd_sc_hd__dfxtp_2
X_786_ _194_ _360_ _361_ _338_ vssd1 vssd1 vccd1 vccd1 _362_ sky130_fd_sc_hd__a31o_1
X_640_ _158_ _171_ _232_ _143_ vssd1 vssd1 vccd1 vccd1 _233_ sky130_fd_sc_hd__a31o_1
X_571_ net15 net35 vssd1 vssd1 vccd1 vccd1 _172_ sky130_fd_sc_hd__and2b_4
X_838_ clknet_3_4__leaf_i_clk _007_ vssd1 vssd1 vccd1 vccd1 o_pc_next[8] sky130_fd_sc_hd__dfxtp_2
X_769_ net26 o_csr_idx[5] _344_ _346_ net23 vssd1 vssd1 vccd1 vccd1 _041_ sky130_fd_sc_hd__o221a_1
X_623_ _170_ _192_ vssd1 vssd1 vccd1 vccd1 _218_ sky130_fd_sc_hd__and2_2
X_554_ i_instruction[0] i_instruction[1] net35 vssd1 vssd1 vccd1 vccd1 _155_ sky130_fd_sc_hd__and3b_1
X_485_ o_funct3[0] _085_ o_funct3[1] vssd1 vssd1 vccd1 vccd1 o_csr_set sky130_fd_sc_hd__and3b_2
X_606_ _158_ _182_ _202_ _146_ vssd1 vssd1 vccd1 vccd1 _203_ sky130_fd_sc_hd__a31o_1
X_537_ _136_ _138_ vssd1 vssd1 vccd1 vccd1 _140_ sky130_fd_sc_hd__nand2_1
X_468_ o_csr_idx[6] net4 net1 vssd1 vssd1 vccd1 vccd1 o_imm_i[26] sky130_fd_sc_hd__a21o_2
X_399_ net40 vssd1 vssd1 vccd1 vccd1 _075_ sky130_fd_sc_hd__inv_2
X_871_ clknet_3_6__leaf_i_clk _040_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[4] sky130_fd_sc_hd__dfxtp_4
X_854_ clknet_3_2__leaf_i_clk _023_ vssd1 vssd1 vccd1 vccd1 o_rd[0] sky130_fd_sc_hd__dfxtp_4
X_785_ _131_ _188_ _340_ _166_ vssd1 vssd1 vccd1 vccd1 _361_ sky130_fd_sc_hd__a211o_1
X_570_ net6 _169_ vssd1 vssd1 vccd1 vccd1 _171_ sky130_fd_sc_hd__nand2_1
X_837_ clknet_3_0__leaf_i_clk _006_ vssd1 vssd1 vccd1 vccd1 o_pc_next[7] sky130_fd_sc_hd__dfxtp_2
X_768_ net12 _345_ net29 vssd1 vssd1 vccd1 vccd1 _346_ sky130_fd_sc_hd__a21o_1
X_699_ _121_ net13 _284_ net31 vssd1 vssd1 vccd1 vccd1 _285_ sky130_fd_sc_hd__a31o_1
X_622_ i_instruction[8] net8 _164_ i_instruction[3] net11 vssd1 vssd1 vccd1 vccd1
+ _217_ sky130_fd_sc_hd__a221o_1
X_553_ _148_ _153_ vssd1 vssd1 vccd1 vccd1 _154_ sky130_fd_sc_hd__nor2_2
X_484_ o_funct3[1] o_funct3[0] _085_ vssd1 vssd1 vccd1 vccd1 o_csr_write sky130_fd_sc_hd__and3b_2
X_605_ i_instruction[6] _173_ vssd1 vssd1 vccd1 vccd1 _202_ sky130_fd_sc_hd__nand2_1
X_536_ _135_ net16 vssd1 vssd1 vccd1 vccd1 _139_ sky130_fd_sc_hd__nor2_2
X_467_ o_csr_idx[5] net4 net1 vssd1 vssd1 vccd1 vccd1 o_imm_i[25] sky130_fd_sc_hd__a21o_2
X_398_ i_instruction[11] vssd1 vssd1 vccd1 vccd1 _074_ sky130_fd_sc_hd__inv_2
Xfanout40 i_instruction[15] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_6
X_519_ net35 i_instruction[10] vssd1 vssd1 vccd1 vccd1 _122_ sky130_fd_sc_hd__and2_2
X_870_ clknet_3_5__leaf_i_clk _039_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[3] sky130_fd_sc_hd__dfxtp_4
X_853_ clknet_3_7__leaf_i_clk _022_ vssd1 vssd1 vccd1 vccd1 instruction\[6\] sky130_fd_sc_hd__dfxtp_4
X_784_ i_instruction[3] _163_ _281_ vssd1 vssd1 vccd1 vccd1 _360_ sky130_fd_sc_hd__a21o_1
X_836_ clknet_3_1__leaf_i_clk _005_ vssd1 vssd1 vccd1 vccd1 o_pc_next[6] sky130_fd_sc_hd__dfxtp_2
X_767_ i_instruction[25] net17 _145_ vssd1 vssd1 vccd1 vccd1 _345_ sky130_fd_sc_hd__mux2_1
X_698_ i_instruction[17] i_instruction[9] _145_ vssd1 vssd1 vccd1 vccd1 _284_ sky130_fd_sc_hd__mux2_1
X_621_ _134_ _151_ vssd1 vssd1 vccd1 vccd1 _216_ sky130_fd_sc_hd__nor2_1
X_552_ i_instruction[5] i_instruction[6] i_instruction[2] i_instruction[3] net36 vssd1
+ vssd1 vccd1 vccd1 _153_ sky130_fd_sc_hd__o41a_1
X_483_ o_csr_idx[5] o_csr_imm_sel _081_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[0] sky130_fd_sc_hd__and3_2
X_819_ o_pc[4] i_pc[4] _114_ vssd1 vssd1 vccd1 vccd1 _051_ sky130_fd_sc_hd__mux2_4
X_604_ net31 instruction\[6\] vssd1 vssd1 vccd1 vccd1 _201_ sky130_fd_sc_hd__nand2_1
X_535_ net33 i_instruction[1] vssd1 vssd1 vccd1 vccd1 _138_ sky130_fd_sc_hd__nand2_4
X_466_ o_csr_idx[4] net4 net1 vssd1 vssd1 vccd1 vccd1 o_imm_i[24] sky130_fd_sc_hd__a21o_2
X_397_ i_instruction[10] vssd1 vssd1 vccd1 vccd1 _073_ sky130_fd_sc_hd__inv_2
Xfanout30 i_stall vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_4
Xfanout41 i_instruction[14] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_6
X_518_ net19 _119_ vssd1 vssd1 vccd1 vccd1 _121_ sky130_fd_sc_hd__or2_4
X_449_ o_rd[0] o_csr_idx[11] _091_ vssd1 vssd1 vccd1 vccd1 _099_ sky130_fd_sc_hd__mux2_1
X_852_ clknet_3_6__leaf_i_clk _021_ vssd1 vssd1 vccd1 vccd1 instruction\[5\] sky130_fd_sc_hd__dfxtp_4
X_783_ net32 _358_ _359_ net25 vssd1 vssd1 vccd1 vccd1 _042_ sky130_fd_sc_hd__o211a_1
X_835_ clknet_3_5__leaf_i_clk _004_ vssd1 vssd1 vccd1 vccd1 o_pc_next[5] sky130_fd_sc_hd__dfxtp_2
X_766_ _338_ _342_ _343_ net11 vssd1 vssd1 vccd1 vccd1 _344_ sky130_fd_sc_hd__o211a_1
X_697_ net5 _282_ _278_ net10 vssd1 vssd1 vccd1 vccd1 _283_ sky130_fd_sc_hd__o211a_1
X_620_ net28 o_rd[0] net25 _215_ vssd1 vssd1 vccd1 vccd1 _023_ sky130_fd_sc_hd__o211a_2
X_551_ _151_ vssd1 vssd1 vccd1 vccd1 _152_ sky130_fd_sc_hd__inv_2
Xclkbuf_3_5__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_482_ _065_ o_funct3[1] _106_ _107_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[2] sky130_fd_sc_hd__a31o_2
X_818_ o_pc[3] i_pc[3] net22 vssd1 vssd1 vccd1 vccd1 _050_ sky130_fd_sc_hd__mux2_2
X_749_ net28 o_csr_idx[3] _323_ _328_ net25 vssd1 vssd1 vccd1 vccd1 _039_ sky130_fd_sc_hd__o221a_2
X_603_ net27 instruction\[5\] net24 _200_ vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__o211a_1
X_534_ net33 i_instruction[1] vssd1 vssd1 vccd1 vccd1 _137_ sky130_fd_sc_hd__and2_2
X_465_ o_csr_idx[3] net4 net1 vssd1 vssd1 vccd1 vccd1 o_imm_i[23] sky130_fd_sc_hd__a21o_2
X_396_ i_instruction[7] vssd1 vssd1 vccd1 vccd1 _072_ sky130_fd_sc_hd__inv_2
Xfanout20 net21 vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_6
Xfanout31 i_stall vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_6
Xfanout42 i_instruction[14] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_4
X_517_ net19 net18 vssd1 vssd1 vccd1 vccd1 _120_ sky130_fd_sc_hd__nor2_4
X_448_ o_alu_ctrl[3] net2 vssd1 vssd1 vccd1 vccd1 o_imm_i[10] sky130_fd_sc_hd__and2_2
X_851_ clknet_3_6__leaf_i_clk _020_ vssd1 vssd1 vccd1 vccd1 instruction\[4\] sky130_fd_sc_hd__dfxtp_2
X_782_ net28 o_csr_idx[6] vssd1 vssd1 vccd1 vccd1 _359_ sky130_fd_sc_hd__or2_1
X_834_ clknet_3_7__leaf_i_clk _003_ vssd1 vssd1 vccd1 vccd1 o_pc_next[4] sky130_fd_sc_hd__dfxtp_2
X_765_ i_instruction[25] _172_ _183_ net17 net7 vssd1 vssd1 vccd1 vccd1 _343_ sky130_fd_sc_hd__a221o_1
X_696_ _218_ _279_ _281_ _257_ vssd1 vssd1 vccd1 vccd1 _282_ sky130_fd_sc_hd__a31o_2
X_550_ net36 i_instruction[3] vssd1 vssd1 vccd1 vccd1 _151_ sky130_fd_sc_hd__nand2_1
X_481_ o_imm_i[10] _104_ _105_ o_inst_branch vssd1 vssd1 vccd1 vccd1 _107_ sky130_fd_sc_hd__a31o_1
X_817_ o_pc[2] i_pc[2] net20 vssd1 vssd1 vccd1 vccd1 _049_ sky130_fd_sc_hd__mux2_1
X_748_ _143_ _326_ _327_ net5 vssd1 vssd1 vccd1 vccd1 _328_ sky130_fd_sc_hd__a22o_1
X_679_ net10 _265_ _266_ _250_ net31 vssd1 vssd1 vccd1 vccd1 _267_ sky130_fd_sc_hd__a221o_1
X_602_ net32 _197_ _198_ _199_ vssd1 vssd1 vccd1 vccd1 _200_ sky130_fd_sc_hd__or4_2
X_533_ net33 i_instruction[0] vssd1 vssd1 vccd1 vccd1 _136_ sky130_fd_sc_hd__nand2_4
X_464_ o_csr_idx[2] net4 net1 vssd1 vssd1 vccd1 vccd1 o_imm_i[22] sky130_fd_sc_hd__a21o_2
X_395_ net39 vssd1 vssd1 vccd1 vccd1 _071_ sky130_fd_sc_hd__inv_2
Xfanout10 net11 vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_4
Xfanout21 _114_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_6
Xfanout32 i_stall vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_4
Xfanout43 i_instruction[13] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_6
X_516_ net34 net40 vssd1 vssd1 vccd1 vccd1 _119_ sky130_fd_sc_hd__and2_4
X_447_ o_csr_idx[9] net3 vssd1 vssd1 vccd1 vccd1 o_imm_i[9] sky130_fd_sc_hd__and2_2
X_850_ clknet_3_7__leaf_i_clk _019_ vssd1 vssd1 vccd1 vccd1 instruction\[3\] sky130_fd_sc_hd__dfxtp_2
X_781_ _353_ _356_ _357_ net10 vssd1 vssd1 vccd1 vccd1 _358_ sky130_fd_sc_hd__o22a_1
X_833_ clknet_3_6__leaf_i_clk _002_ vssd1 vssd1 vccd1 vccd1 o_pc_next[3] sky130_fd_sc_hd__dfxtp_2
X_764_ _281_ _339_ _341_ _194_ vssd1 vssd1 vccd1 vccd1 _342_ sky130_fd_sc_hd__o211a_1
X_695_ _166_ _280_ vssd1 vssd1 vccd1 vccd1 _281_ sky130_fd_sc_hd__nand2_2
X_480_ o_csr_idx[5] instruction\[6\] _080_ _105_ vssd1 vssd1 vccd1 vccd1 _106_ sky130_fd_sc_hd__o31ai_1
X_816_ o_pc[1] i_pc[1] net20 vssd1 vssd1 vccd1 vccd1 _048_ sky130_fd_sc_hd__mux2_1
X_747_ i_instruction[23] _135_ net15 net39 vssd1 vssd1 vccd1 vccd1 _327_ sky130_fd_sc_hd__a22o_1
X_678_ _072_ net19 vssd1 vssd1 vccd1 vccd1 _266_ sky130_fd_sc_hd__nand2_1
X_601_ net39 _135_ net16 _156_ vssd1 vssd1 vccd1 vccd1 _199_ sky130_fd_sc_hd__a31o_1
X_532_ net35 i_instruction[0] vssd1 vssd1 vccd1 vccd1 _135_ sky130_fd_sc_hd__and2_4
X_463_ o_csr_idx[1] net4 net1 vssd1 vssd1 vccd1 vccd1 o_imm_i[21] sky130_fd_sc_hd__a21o_2
X_394_ i_flush vssd1 vssd1 vccd1 vccd1 _070_ sky130_fd_sc_hd__inv_2
Xfanout11 _140_ vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_4
Xfanout22 _114_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_12
Xfanout33 net38 vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_8
X_515_ net33 net41 vssd1 vssd1 vccd1 vccd1 _118_ sky130_fd_sc_hd__nand2_8
X_446_ o_csr_idx[8] net2 vssd1 vssd1 vccd1 vccd1 o_imm_i[8] sky130_fd_sc_hd__and2_2
X_429_ _090_ vssd1 vssd1 vccd1 vccd1 o_inst_store sky130_fd_sc_hd__inv_2
X_780_ net39 _117_ net9 i_instruction[26] _262_ vssd1 vssd1 vccd1 vccd1 _357_ sky130_fd_sc_hd__a221o_1
X_901_ o_csr_idx[4] vssd1 vssd1 vccd1 vccd1 o_rs2[4] sky130_fd_sc_hd__buf_2
X_832_ clknet_3_1__leaf_i_clk _001_ vssd1 vssd1 vccd1 vccd1 o_pc_next[2] sky130_fd_sc_hd__dfxtp_2
X_763_ net34 i_instruction[2] _188_ _340_ _166_ vssd1 vssd1 vccd1 vccd1 _341_ sky130_fd_sc_hd__a311o_1
X_694_ _124_ _162_ _130_ vssd1 vssd1 vccd1 vccd1 _280_ sky130_fd_sc_hd__a21o_1
X_815_ net23 _386_ vssd1 vssd1 vccd1 vccd1 _047_ sky130_fd_sc_hd__and2_1
X_746_ net34 net39 _120_ _325_ vssd1 vssd1 vccd1 vccd1 _326_ sky130_fd_sc_hd__a31o_1
X_677_ _138_ _260_ _264_ _160_ vssd1 vssd1 vccd1 vccd1 _265_ sky130_fd_sc_hd__a22o_1
X_600_ i_instruction[5] net19 net18 net12 vssd1 vssd1 vccd1 vccd1 _198_ sky130_fd_sc_hd__o211a_1
X_531_ _128_ _130_ _132_ _121_ vssd1 vssd1 vccd1 vccd1 _134_ sky130_fd_sc_hd__a31o_1
X_462_ o_csr_idx[0] _088_ _101_ vssd1 vssd1 vccd1 vccd1 o_imm_i[20] sky130_fd_sc_hd__a21o_2
X_393_ instruction\[2\] vssd1 vssd1 vccd1 vccd1 _069_ sky130_fd_sc_hd__inv_2
X_729_ net11 _310_ vssd1 vssd1 vccd1 vccd1 _311_ sky130_fd_sc_hd__and2_1
Xfanout12 _139_ vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_6
Xfanout23 net25 vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_4
Xfanout34 net35 vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_4
X_514_ net33 net41 vssd1 vssd1 vccd1 vccd1 _117_ sky130_fd_sc_hd__and2_2
X_445_ o_csr_idx[7] net3 vssd1 vssd1 vccd1 vccd1 o_imm_i[7] sky130_fd_sc_hd__and2_2
X_428_ instruction\[5\] _083_ vssd1 vssd1 vccd1 vccd1 _090_ sky130_fd_sc_hd__nand2_1
X_900_ o_csr_idx[3] vssd1 vssd1 vccd1 vccd1 o_rs2[3] sky130_fd_sc_hd__buf_2
X_831_ clknet_3_0__leaf_i_clk _000_ vssd1 vssd1 vccd1 vccd1 o_pc_next[1] sky130_fd_sc_hd__dfxtp_2
X_762_ _073_ i_instruction[12] _123_ _187_ vssd1 vssd1 vccd1 vccd1 _340_ sky130_fd_sc_hd__and4_2
X_693_ net36 i_instruction[9] _166_ vssd1 vssd1 vccd1 vccd1 _279_ sky130_fd_sc_hd__a21o_1
X_814_ o_csr_idx[11] net29 _147_ _385_ vssd1 vssd1 vccd1 vccd1 _386_ sky130_fd_sc_hd__a22o_1
X_745_ i_instruction[10] net19 net18 _324_ net30 vssd1 vssd1 vccd1 vccd1 _325_ sky130_fd_sc_hd__a221o_1
X_676_ net18 net14 _261_ _263_ vssd1 vssd1 vccd1 vccd1 _264_ sky130_fd_sc_hd__o22a_1
X_530_ _128_ _130_ _132_ _121_ vssd1 vssd1 vccd1 vccd1 _133_ sky130_fd_sc_hd__a31oi_4
X_461_ o_csr_imm[4] _094_ _102_ vssd1 vssd1 vccd1 vccd1 o_imm_i[19] sky130_fd_sc_hd__a21o_2
X_392_ instruction\[3\] vssd1 vssd1 vccd1 vccd1 _068_ sky130_fd_sc_hd__inv_2
X_728_ i_instruction[21] _173_ _308_ net7 _309_ vssd1 vssd1 vccd1 vccd1 _310_ sky130_fd_sc_hd__a221o_1
X_659_ _169_ _247_ _248_ _240_ vssd1 vssd1 vccd1 vccd1 _249_ sky130_fd_sc_hd__o31a_1
Xfanout13 _139_ vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_2
Xfanout24 net25 vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_2
Xfanout35 net37 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_8
X_513_ net31 instruction\[0\] vssd1 vssd1 vccd1 vccd1 _116_ sky130_fd_sc_hd__nand2_1
X_444_ o_csr_idx[6] net3 vssd1 vssd1 vccd1 vccd1 o_imm_i[6] sky130_fd_sc_hd__and2_2
X_427_ o_csr_imm[4] net2 vssd1 vssd1 vccd1 vccd1 o_rs1[4] sky130_fd_sc_hd__and2_2
X_830_ o_pc[15] i_pc[15] net20 vssd1 vssd1 vccd1 vccd1 _062_ sky130_fd_sc_hd__mux2_1
X_761_ i_instruction[2] _124_ _162_ vssd1 vssd1 vccd1 vccd1 _339_ sky130_fd_sc_hd__and3_1
X_692_ i_instruction[9] net14 _276_ _277_ vssd1 vssd1 vccd1 vccd1 _278_ sky130_fd_sc_hd__a31o_1
X_813_ i_instruction[31] _173_ _369_ net7 vssd1 vssd1 vccd1 vccd1 _385_ sky130_fd_sc_hd__a22o_1
X_744_ net42 i_instruction[23] vssd1 vssd1 vccd1 vccd1 _324_ sky130_fd_sc_hd__or2_1
X_675_ _121_ _125_ net14 vssd1 vssd1 vccd1 vccd1 _263_ sky130_fd_sc_hd__o21ai_1
X_460_ o_csr_imm[3] _094_ _102_ vssd1 vssd1 vccd1 vccd1 o_imm_i[18] sky130_fd_sc_hd__a21o_2
X_391_ instruction\[4\] vssd1 vssd1 vccd1 vccd1 _067_ sky130_fd_sc_hd__clkinv_2
X_727_ i_instruction[3] net15 _165_ vssd1 vssd1 vccd1 vccd1 _309_ sky130_fd_sc_hd__and3_1
X_658_ i_instruction[6] _073_ _123_ _187_ vssd1 vssd1 vccd1 vccd1 _248_ sky130_fd_sc_hd__o211a_1
X_589_ net42 i_instruction[13] net40 net34 vssd1 vssd1 vccd1 vccd1 _187_ sky130_fd_sc_hd__and4bb_4
Xfanout14 net15 vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_4
Xfanout25 _070_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_6
Xfanout36 net37 vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_6
X_512_ net27 valid_input net24 _115_ vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__o211a_1
X_443_ o_csr_idx[5] net3 vssd1 vssd1 vccd1 vccd1 o_imm_i[5] sky130_fd_sc_hd__and2_2
X_426_ o_csr_imm[3] net3 vssd1 vssd1 vccd1 vccd1 o_rs1[3] sky130_fd_sc_hd__and2_2
X_409_ instruction\[6\] _080_ vssd1 vssd1 vccd1 vccd1 _081_ sky130_fd_sc_hd__nor2_2
X_760_ net17 _193_ net5 vssd1 vssd1 vccd1 vccd1 _338_ sky130_fd_sc_hd__a21o_1
X_691_ i_instruction[17] _172_ net6 vssd1 vssd1 vccd1 vccd1 _277_ sky130_fd_sc_hd__a21o_1
X_889_ clknet_3_4__leaf_i_clk _058_ vssd1 vssd1 vccd1 vccd1 o_pc[11] sky130_fd_sc_hd__dfxtp_2
X_812_ _070_ _384_ vssd1 vssd1 vccd1 vccd1 _046_ sky130_fd_sc_hd__and2_1
X_743_ _293_ _321_ _322_ net7 vssd1 vssd1 vccd1 vccd1 _323_ sky130_fd_sc_hd__o31a_1
X_674_ _121_ _125_ vssd1 vssd1 vccd1 vccd1 _262_ sky130_fd_sc_hd__nor2_1
X_390_ instruction\[6\] vssd1 vssd1 vccd1 vccd1 _066_ sky130_fd_sc_hd__inv_2
X_726_ _152_ _307_ _293_ vssd1 vssd1 vccd1 vccd1 _308_ sky130_fd_sc_hd__a21o_1
X_657_ _151_ _168_ vssd1 vssd1 vccd1 vccd1 _247_ sky130_fd_sc_hd__nor2_1
X_588_ net27 instruction\[4\] net24 _186_ vssd1 vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__o211a_1
Xfanout15 _155_ vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_4
Xfanout26 net28 vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_4
Xfanout37 net38 vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_4
X_511_ net29 net38 vssd1 vssd1 vccd1 vccd1 _115_ sky130_fd_sc_hd__or2_1
X_442_ net2 _098_ vssd1 vssd1 vccd1 vccd1 o_imm_i[4] sky130_fd_sc_hd__and2_2
X_709_ _130_ _168_ vssd1 vssd1 vccd1 vccd1 _293_ sky130_fd_sc_hd__nor2_4
X_425_ o_csr_imm[2] net3 vssd1 vssd1 vccd1 vccd1 o_rs1[2] sky130_fd_sc_hd__and2_2
X_408_ instruction\[5\] instruction\[4\] _076_ vssd1 vssd1 vccd1 vccd1 _080_ sky130_fd_sc_hd__nand3_2
X_690_ net19 _268_ vssd1 vssd1 vccd1 vccd1 _276_ sky130_fd_sc_hd__nor2_1
X_888_ clknet_3_2__leaf_i_clk _057_ vssd1 vssd1 vccd1 vccd1 o_pc[10] sky130_fd_sc_hd__dfxtp_2
X_811_ net30 o_alu_ctrl[3] _147_ _383_ vssd1 vssd1 vccd1 vccd1 _384_ sky130_fd_sc_hd__a22o_1
X_742_ net35 _073_ _074_ _188_ vssd1 vssd1 vccd1 vccd1 _322_ sky130_fd_sc_hd__a211oi_1
X_673_ net17 _154_ net8 i_instruction[7] vssd1 vssd1 vccd1 vccd1 _261_ sky130_fd_sc_hd__o211a_1
Xclkbuf_3_1__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_725_ net42 _194_ vssd1 vssd1 vccd1 vccd1 _307_ sky130_fd_sc_hd__nand2_1
X_656_ net23 _246_ vssd1 vssd1 vccd1 vccd1 _028_ sky130_fd_sc_hd__and2_1
X_587_ _180_ _182_ _185_ net32 vssd1 vssd1 vccd1 vccd1 _186_ sky130_fd_sc_hd__a31o_1
Xfanout16 _137_ vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_6
Xfanout27 net28 vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_4
Xfanout38 i_ready vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_4
X_510_ o_pc_next[15] i_pc_next[15] net21 vssd1 vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__mux2_1
X_441_ o_rd[4] o_csr_idx[4] _092_ vssd1 vssd1 vccd1 vccd1 _098_ sky130_fd_sc_hd__mux2_1
X_708_ i_instruction[19] _172_ _291_ net7 vssd1 vssd1 vccd1 vccd1 _292_ sky130_fd_sc_hd__a211o_1
X_639_ net9 net6 _122_ vssd1 vssd1 vccd1 vccd1 _232_ sky130_fd_sc_hd__a21o_1
X_424_ o_csr_imm[1] net2 vssd1 vssd1 vccd1 vccd1 o_rs1[1] sky130_fd_sc_hd__and2_2
X_407_ _068_ _078_ vssd1 vssd1 vccd1 vccd1 o_inst_jal sky130_fd_sc_hd__nor2_4
X_887_ clknet_3_5__leaf_i_clk _056_ vssd1 vssd1 vccd1 vccd1 o_pc[9] sky130_fd_sc_hd__dfxtp_2
X_810_ i_instruction[30] _173_ _382_ net7 vssd1 vssd1 vccd1 vccd1 _383_ sky130_fd_sc_hd__a22o_1
X_741_ net34 net39 _307_ vssd1 vssd1 vccd1 vccd1 _321_ sky130_fd_sc_hd__and3_1
X_672_ _218_ _258_ _259_ _257_ vssd1 vssd1 vccd1 vccd1 _260_ sky130_fd_sc_hd__a31o_1
X_724_ net26 o_csr_idx[0] net23 _306_ vssd1 vssd1 vccd1 vccd1 _036_ sky130_fd_sc_hd__o211a_1
X_655_ net29 o_funct3[0] _147_ _245_ vssd1 vssd1 vccd1 vccd1 _246_ sky130_fd_sc_hd__a22o_1
X_586_ _179_ _183_ _184_ _137_ vssd1 vssd1 vccd1 vccd1 _185_ sky130_fd_sc_hd__o31ai_1
Xfanout17 _129_ vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_4
Xfanout28 _063_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_6
Xfanout39 i_instruction[5] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_6
X_440_ net2 _097_ vssd1 vssd1 vccd1 vccd1 o_imm_i[3] sky130_fd_sc_hd__and2_2
X_707_ net41 _268_ net15 i_instruction[11] vssd1 vssd1 vccd1 vccd1 _291_ sky130_fd_sc_hd__and4bb_1
X_638_ net27 o_rd[2] net24 _231_ vssd1 vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__o211a_1
X_569_ net35 net43 _118_ vssd1 vssd1 vccd1 vccd1 _170_ sky130_fd_sc_hd__nand3_4
X_423_ o_csr_imm[0] net3 vssd1 vssd1 vccd1 vccd1 o_rs1[0] sky130_fd_sc_hd__and2_2
X_406_ instruction\[3\] _077_ vssd1 vssd1 vccd1 vccd1 _079_ sky130_fd_sc_hd__and2_1
X_886_ clknet_3_1__leaf_i_clk _055_ vssd1 vssd1 vccd1 vccd1 o_pc[8] sky130_fd_sc_hd__dfxtp_2
X_740_ net26 o_csr_idx[2] net23 _320_ vssd1 vssd1 vccd1 vccd1 _038_ sky130_fd_sc_hd__o211a_1
X_671_ _125_ _165_ vssd1 vssd1 vccd1 vccd1 _259_ sky130_fd_sc_hd__nand2_1
X_869_ clknet_3_4__leaf_i_clk _038_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[2] sky130_fd_sc_hd__dfxtp_4
X_723_ net16 _301_ _303_ _305_ vssd1 vssd1 vccd1 vccd1 _306_ sky130_fd_sc_hd__a211o_1
X_654_ _239_ _240_ _242_ _244_ vssd1 vssd1 vccd1 vccd1 _245_ sky130_fd_sc_hd__a31o_1
X_585_ _148_ net14 vssd1 vssd1 vccd1 vccd1 _184_ sky130_fd_sc_hd__nor2_1
Xfanout18 _119_ vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_6
Xfanout29 i_stall vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_6
X_706_ net26 o_csr_imm[3] _288_ _290_ net23 vssd1 vssd1 vccd1 vccd1 _034_ sky130_fd_sc_hd__o221a_1
X_637_ _227_ _228_ _230_ net32 vssd1 vssd1 vccd1 vccd1 _231_ sky130_fd_sc_hd__a31o_1
X_568_ net33 net43 _118_ vssd1 vssd1 vccd1 vccd1 _169_ sky130_fd_sc_hd__and3_4
X_499_ o_pc_next[4] i_pc_next[4] net22 vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__mux2_2
X_422_ _067_ instruction\[3\] _069_ vssd1 vssd1 vccd1 vccd1 _089_ sky130_fd_sc_hd__or3_2
X_405_ instruction\[3\] _078_ vssd1 vssd1 vccd1 vccd1 o_inst_jalr sky130_fd_sc_hd__nor2_4
X_885_ clknet_3_1__leaf_i_clk _054_ vssd1 vssd1 vccd1 vccd1 o_pc[7] sky130_fd_sc_hd__dfxtp_2
X_670_ _071_ _163_ _164_ vssd1 vssd1 vccd1 vccd1 _258_ sky130_fd_sc_hd__o21ai_1
X_868_ clknet_3_1__leaf_i_clk _037_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[1] sky130_fd_sc_hd__dfxtp_4
X_799_ i_instruction[28] _138_ _135_ vssd1 vssd1 vccd1 vccd1 _374_ sky130_fd_sc_hd__o21a_1
X_722_ _257_ _293_ _304_ net7 vssd1 vssd1 vccd1 vccd1 _305_ sky130_fd_sc_hd__o31a_1
X_653_ net17 net14 net5 _243_ vssd1 vssd1 vccd1 vccd1 _244_ sky130_fd_sc_hd__o211a_1
X_584_ net41 net15 vssd1 vssd1 vccd1 vccd1 _183_ sky130_fd_sc_hd__and2_1
Xfanout19 _117_ vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_6
X_705_ net16 _286_ _289_ _250_ net29 vssd1 vssd1 vccd1 vccd1 _290_ sky130_fd_sc_hd__a221o_1
X_636_ net38 i_instruction[9] _182_ _229_ vssd1 vssd1 vccd1 vccd1 _230_ sky130_fd_sc_hd__a31o_1
X_567_ _124_ _162_ _167_ vssd1 vssd1 vccd1 vccd1 _168_ sky130_fd_sc_hd__a21o_4
X_498_ o_pc_next[3] i_pc_next[3] net22 vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__mux2_2
X_421_ instruction\[4\] _068_ instruction\[2\] vssd1 vssd1 vccd1 vccd1 _088_ sky130_fd_sc_hd__and3_4
X_619_ _208_ _212_ _214_ net32 vssd1 vssd1 vccd1 vccd1 _215_ sky130_fd_sc_hd__a31o_1
X_404_ _078_ vssd1 vssd1 vccd1 vccd1 o_res_src[1] sky130_fd_sc_hd__clkinv_4
Xclkbuf_3_4__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_884_ clknet_3_5__leaf_i_clk _053_ vssd1 vssd1 vccd1 vccd1 o_pc[6] sky130_fd_sc_hd__dfxtp_2
X_867_ clknet_3_5__leaf_i_clk _036_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[0] sky130_fd_sc_hd__dfxtp_4
X_798_ _371_ _372_ net16 vssd1 vssd1 vccd1 vccd1 _373_ sky130_fd_sc_hd__a21o_1
X_721_ _188_ _194_ _150_ vssd1 vssd1 vccd1 vccd1 _304_ sky130_fd_sc_hd__a21oi_1
X_652_ _121_ net15 vssd1 vssd1 vccd1 vccd1 _243_ sky130_fd_sc_hd__nand2_1
X_583_ net6 _181_ vssd1 vssd1 vccd1 vccd1 _182_ sky130_fd_sc_hd__nand2_1
X_704_ i_instruction[18] _117_ vssd1 vssd1 vccd1 vccd1 _289_ sky130_fd_sc_hd__or2_1
X_635_ i_instruction[15] i_instruction[4] net19 net13 vssd1 vssd1 vccd1 vccd1 _229_
+ sky130_fd_sc_hd__a31o_1
X_566_ net40 net43 net36 net42 vssd1 vssd1 vccd1 vccd1 _167_ sky130_fd_sc_hd__nand4b_1
X_497_ o_pc_next[2] i_pc_next[2] net20 vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__mux2_1
X_420_ o_csr_idx[2] _064_ _086_ o_csr_idx[9] vssd1 vssd1 vccd1 vccd1 o_inst_mret sky130_fd_sc_hd__nor4b_4
X_618_ net36 i_instruction[2] _133_ _213_ vssd1 vssd1 vccd1 vccd1 _214_ sky130_fd_sc_hd__a31o_1
X_549_ net36 i_instruction[2] vssd1 vssd1 vccd1 vccd1 _150_ sky130_fd_sc_hd__nand2_2
X_403_ instruction\[2\] _077_ vssd1 vssd1 vccd1 vccd1 _078_ sky130_fd_sc_hd__nand2_8
X_883_ clknet_3_0__leaf_i_clk _052_ vssd1 vssd1 vccd1 vccd1 o_pc[5] sky130_fd_sc_hd__dfxtp_2
X_866_ clknet_3_3__leaf_i_clk _035_ vssd1 vssd1 vccd1 vccd1 o_csr_imm[4] sky130_fd_sc_hd__dfxtp_4
X_797_ i_instruction[9] _170_ _370_ _166_ vssd1 vssd1 vccd1 vccd1 _372_ sky130_fd_sc_hd__o22a_1
X_720_ net18 net12 _302_ net30 vssd1 vssd1 vccd1 vccd1 _303_ sky130_fd_sc_hd__a31o_1
X_651_ _150_ _163_ _166_ vssd1 vssd1 vccd1 vccd1 _242_ sky130_fd_sc_hd__o21ai_1
X_582_ net41 net43 _165_ net38 vssd1 vssd1 vccd1 vccd1 _181_ sky130_fd_sc_hd__o211a_1
X_849_ clknet_3_3__leaf_i_clk _018_ vssd1 vssd1 vccd1 vccd1 instruction\[2\] sky130_fd_sc_hd__dfxtp_4
X_703_ i_instruction[10] _196_ _287_ net6 vssd1 vssd1 vccd1 vccd1 _288_ sky130_fd_sc_hd__o211a_1
X_634_ i_instruction[9] _158_ _138_ vssd1 vssd1 vccd1 vccd1 _228_ sky130_fd_sc_hd__a21o_1
X_565_ net40 i_instruction[13] net34 net42 vssd1 vssd1 vccd1 vccd1 _166_ sky130_fd_sc_hd__and4b_4
X_496_ o_pc_next[1] i_pc_next[1] net21 vssd1 vssd1 vccd1 vccd1 _000_ sky130_fd_sc_hd__mux2_1
X_617_ i_instruction[7] net9 _164_ i_instruction[2] net11 vssd1 vssd1 vccd1 vccd1
+ _213_ sky130_fd_sc_hd__a221o_1
X_548_ net33 i_instruction[4] vssd1 vssd1 vccd1 vccd1 _149_ sky130_fd_sc_hd__nand2_1
X_479_ instruction\[2\] _103_ vssd1 vssd1 vccd1 vccd1 _105_ sky130_fd_sc_hd__or2_1
X_402_ _076_ _077_ vssd1 vssd1 vccd1 vccd1 o_inst_branch sky130_fd_sc_hd__and2_4
X_882_ clknet_3_5__leaf_i_clk _051_ vssd1 vssd1 vccd1 vccd1 o_pc[4] sky130_fd_sc_hd__dfxtp_2
X_865_ clknet_3_7__leaf_i_clk _034_ vssd1 vssd1 vccd1 vccd1 o_csr_imm[3] sky130_fd_sc_hd__dfxtp_4
X_796_ _148_ _163_ _281_ vssd1 vssd1 vccd1 vccd1 _371_ sky130_fd_sc_hd__a21o_1
X_650_ _240_ vssd1 vssd1 vccd1 vccd1 _241_ sky130_fd_sc_hd__inv_2
X_581_ i_instruction[4] net9 net10 _133_ vssd1 vssd1 vccd1 vccd1 _180_ sky130_fd_sc_hd__a211o_1
X_848_ clknet_3_6__leaf_i_clk _017_ vssd1 vssd1 vccd1 vccd1 instruction\[1\] sky130_fd_sc_hd__dfxtp_1
X_779_ i_instruction[1] _355_ net13 vssd1 vssd1 vccd1 vccd1 _356_ sky130_fd_sc_hd__a21o_1
X_702_ _218_ _281_ _257_ vssd1 vssd1 vccd1 vccd1 _287_ sky130_fd_sc_hd__a21o_1
X_633_ _148_ _225_ _226_ net10 vssd1 vssd1 vccd1 vccd1 _227_ sky130_fd_sc_hd__a211o_1
X_564_ net40 net42 net34 vssd1 vssd1 vccd1 vccd1 _165_ sky130_fd_sc_hd__nand3b_4
X_495_ net31 i_flush vssd1 vssd1 vccd1 vccd1 _114_ sky130_fd_sc_hd__nor2_8
X_616_ _128_ _145_ _210_ _211_ vssd1 vssd1 vccd1 vccd1 _212_ sky130_fd_sc_hd__o31ai_1
X_547_ net35 i_instruction[4] vssd1 vssd1 vccd1 vccd1 _148_ sky130_fd_sc_hd__and2_4
X_478_ net2 _104_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[4] sky130_fd_sc_hd__nand2_4
X_401_ instruction\[6\] instruction\[5\] _067_ vssd1 vssd1 vccd1 vccd1 _077_ sky130_fd_sc_hd__and3_2
X_881_ clknet_3_7__leaf_i_clk _050_ vssd1 vssd1 vccd1 vccd1 o_pc[3] sky130_fd_sc_hd__dfxtp_2
X_864_ clknet_3_2__leaf_i_clk _033_ vssd1 vssd1 vccd1 vccd1 o_csr_imm[2] sky130_fd_sc_hd__dfxtp_4
X_795_ net17 _188_ _340_ _169_ vssd1 vssd1 vccd1 vccd1 _370_ sky130_fd_sc_hd__a211o_1
X_580_ _161_ _157_ vssd1 vssd1 vccd1 vccd1 _179_ sky130_fd_sc_hd__and2b_1
X_847_ clknet_3_3__leaf_i_clk _016_ vssd1 vssd1 vccd1 vccd1 instruction\[0\] sky130_fd_sc_hd__dfxtp_1
X_778_ i_instruction[26] _135_ _259_ _354_ vssd1 vssd1 vccd1 vccd1 _355_ sky130_fd_sc_hd__a22o_1
X_701_ i_instruction[10] _136_ _276_ _172_ i_instruction[18] vssd1 vssd1 vccd1 vccd1
+ _286_ sky130_fd_sc_hd__a32o_1
X_632_ i_instruction[9] net41 _118_ i_instruction[6] _119_ vssd1 vssd1 vccd1 vccd1
+ _226_ sky130_fd_sc_hd__o221a_1
X_563_ i_instruction[15] net42 net37 vssd1 vssd1 vccd1 vccd1 _164_ sky130_fd_sc_hd__and3b_2
X_494_ _087_ o_inst_mret _111_ _113_ vssd1 vssd1 vccd1 vccd1 o_inst_supported sky130_fd_sc_hd__or4b_4
Xclkbuf_3_7__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_615_ _072_ net16 _156_ vssd1 vssd1 vccd1 vccd1 _211_ sky130_fd_sc_hd__a21o_1
X_546_ net12 _145_ net29 vssd1 vssd1 vccd1 vccd1 _147_ sky130_fd_sc_hd__a21oi_4
X_477_ o_inst_jal _083_ vssd1 vssd1 vccd1 vccd1 _104_ sky130_fd_sc_hd__nor2_4
X_400_ instruction\[3\] instruction\[2\] vssd1 vssd1 vccd1 vccd1 _076_ sky130_fd_sc_hd__nor2_2
X_529_ net39 i_instruction[6] net35 vssd1 vssd1 vccd1 vccd1 _132_ sky130_fd_sc_hd__o21ai_4
X_880_ clknet_3_4__leaf_i_clk _049_ vssd1 vssd1 vccd1 vccd1 o_pc[2] sky130_fd_sc_hd__dfxtp_2
X_863_ clknet_3_3__leaf_i_clk _032_ vssd1 vssd1 vccd1 vccd1 o_csr_imm[1] sky130_fd_sc_hd__dfxtp_4
X_794_ net17 _188_ _340_ vssd1 vssd1 vccd1 vccd1 _369_ sky130_fd_sc_hd__a21o_1
X_846_ clknet_3_6__leaf_i_clk _015_ vssd1 vssd1 vccd1 vccd1 valid_input sky130_fd_sc_hd__dfxtp_1
X_777_ i_instruction[2] net18 net14 net19 vssd1 vssd1 vccd1 vccd1 _354_ sky130_fd_sc_hd__o211a_1
X_700_ net27 o_csr_imm[2] _283_ _285_ net24 vssd1 vssd1 vccd1 vccd1 _033_ sky130_fd_sc_hd__o221a_2
X_631_ _134_ _165_ vssd1 vssd1 vccd1 vccd1 _225_ sky130_fd_sc_hd__nand2_1
X_562_ _124_ _162_ vssd1 vssd1 vccd1 vccd1 _163_ sky130_fd_sc_hd__and2_2
X_493_ _078_ _084_ _112_ _091_ valid_input vssd1 vssd1 vccd1 vccd1 _113_ sky130_fd_sc_hd__o311a_1
X_829_ o_pc[14] i_pc[14] net21 vssd1 vssd1 vccd1 vccd1 _061_ sky130_fd_sc_hd__mux2_1
X_614_ _125_ _154_ _209_ vssd1 vssd1 vccd1 vccd1 _210_ sky130_fd_sc_hd__o21ba_1
X_545_ _136_ _138_ _145_ net30 vssd1 vssd1 vccd1 vccd1 _146_ sky130_fd_sc_hd__a31o_1
X_476_ o_csr_idx[5] _081_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[1] sky130_fd_sc_hd__and2_2
X_528_ net37 i_instruction[6] vssd1 vssd1 vccd1 vccd1 _131_ sky130_fd_sc_hd__and2_2
X_459_ o_csr_imm[2] _094_ _102_ vssd1 vssd1 vccd1 vccd1 o_imm_i[17] sky130_fd_sc_hd__a21o_2
X_862_ clknet_3_6__leaf_i_clk _031_ vssd1 vssd1 vccd1 vccd1 o_csr_imm[0] sky130_fd_sc_hd__dfxtp_4
X_793_ _143_ _366_ _368_ net32 _367_ vssd1 vssd1 vccd1 vccd1 _043_ sky130_fd_sc_hd__o221a_2
X_845_ clknet_3_0__leaf_i_clk _014_ vssd1 vssd1 vccd1 vccd1 o_pc_next[15] sky130_fd_sc_hd__dfxtp_2
X_776_ _196_ _351_ _352_ vssd1 vssd1 vccd1 vccd1 _353_ sky130_fd_sc_hd__a21oi_1
X_630_ net31 _223_ _224_ net24 vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__o211a_2
X_561_ i_instruction[7] i_instruction[8] net37 vssd1 vssd1 vccd1 vccd1 _162_ sky130_fd_sc_hd__and3b_1
X_492_ o_csr_imm_sel o_funct3[1] o_funct3[0] _068_ vssd1 vssd1 vccd1 vccd1 _112_ sky130_fd_sc_hd__o31a_1
X_828_ o_pc[13] i_pc[13] net22 vssd1 vssd1 vccd1 vccd1 _060_ sky130_fd_sc_hd__mux2_1
X_759_ _063_ o_csr_idx[4] _336_ _337_ _070_ vssd1 vssd1 vccd1 vccd1 _040_ sky130_fd_sc_hd__o221a_1
X_613_ net17 _154_ net14 _165_ vssd1 vssd1 vccd1 vccd1 _209_ sky130_fd_sc_hd__and4_1
X_544_ net41 net40 net33 vssd1 vssd1 vccd1 vccd1 _145_ sky130_fd_sc_hd__nand3b_4
X_475_ _069_ _103_ o_inst_jal vssd1 vssd1 vccd1 vccd1 o_op1_src sky130_fd_sc_hd__o21bai_4
X_527_ net36 i_instruction[12] vssd1 vssd1 vccd1 vccd1 _130_ sky130_fd_sc_hd__nand2_8
X_458_ o_csr_imm[1] _094_ _102_ vssd1 vssd1 vccd1 vccd1 o_imm_i[16] sky130_fd_sc_hd__a21o_2
X_389_ o_csr_imm_sel vssd1 vssd1 vccd1 vccd1 _065_ sky130_fd_sc_hd__inv_2
X_861_ clknet_3_7__leaf_i_clk _030_ vssd1 vssd1 vccd1 vccd1 o_csr_imm_sel sky130_fd_sc_hd__dfxtp_4
X_792_ _120_ _126_ net8 i_instruction[27] net10 vssd1 vssd1 vccd1 vccd1 _368_ sky130_fd_sc_hd__a221o_1
X_844_ clknet_3_5__leaf_i_clk _013_ vssd1 vssd1 vccd1 vccd1 o_pc_next[14] sky130_fd_sc_hd__dfxtp_2
X_775_ _130_ _193_ _160_ vssd1 vssd1 vccd1 vccd1 _352_ sky130_fd_sc_hd__a21o_1
X_560_ _128_ net17 vssd1 vssd1 vccd1 vccd1 _161_ sky130_fd_sc_hd__and2_1
X_491_ _084_ _110_ o_csr_read vssd1 vssd1 vccd1 vccd1 _111_ sky130_fd_sc_hd__o21bai_1
X_827_ o_pc[12] i_pc[12] net21 vssd1 vssd1 vccd1 vccd1 _059_ sky130_fd_sc_hd__mux2_1
X_758_ net6 _196_ _329_ _333_ vssd1 vssd1 vccd1 vccd1 _337_ sky130_fd_sc_hd__a31o_1
X_689_ net28 o_csr_imm[1] _273_ _275_ net25 vssd1 vssd1 vccd1 vccd1 _032_ sky130_fd_sc_hd__o221a_2
X_612_ i_instruction[7] _195_ _207_ net5 vssd1 vssd1 vccd1 vccd1 _208_ sky130_fd_sc_hd__a211o_1
X_543_ _118_ net18 vssd1 vssd1 vccd1 vccd1 _144_ sky130_fd_sc_hd__and2_1
X_474_ instruction\[6\] instruction\[5\] _067_ instruction\[3\] vssd1 vssd1 vccd1
+ vccd1 _103_ sky130_fd_sc_hd__or4_2
X_526_ net37 i_instruction[12] vssd1 vssd1 vccd1 vccd1 _129_ sky130_fd_sc_hd__and2_1
X_457_ o_csr_imm[0] _094_ _102_ vssd1 vssd1 vccd1 vccd1 o_imm_i[15] sky130_fd_sc_hd__a21o_2
X_388_ o_csr_idx[1] vssd1 vssd1 vccd1 vccd1 _064_ sky130_fd_sc_hd__clkinv_2
Xclkbuf_3_0__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_509_ o_pc_next[14] i_pc_next[14] net22 vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__mux2_2
X_860_ clknet_3_4__leaf_i_clk _029_ vssd1 vssd1 vccd1 vccd1 o_funct3[1] sky130_fd_sc_hd__dfxtp_4
X_791_ net28 o_csr_idx[7] net25 vssd1 vssd1 vccd1 vccd1 _367_ sky130_fd_sc_hd__o21a_1
X_843_ clknet_3_3__leaf_i_clk _012_ vssd1 vssd1 vccd1 vccd1 o_pc_next[13] sky130_fd_sc_hd__dfxtp_2
X_774_ _218_ _348_ _350_ _169_ _072_ vssd1 vssd1 vccd1 vccd1 _351_ sky130_fd_sc_hd__a32o_1
X_490_ instruction\[4\] _068_ _069_ _108_ _109_ vssd1 vssd1 vccd1 vccd1 _110_ sky130_fd_sc_hd__o41a_1
X_826_ o_pc[11] i_pc[11] net20 vssd1 vssd1 vccd1 vccd1 _058_ sky130_fd_sc_hd__mux2_1
X_757_ i_instruction[6] net6 _335_ vssd1 vssd1 vccd1 vccd1 _336_ sky130_fd_sc_hd__and3_1
X_688_ net31 _133_ _274_ _143_ vssd1 vssd1 vccd1 vccd1 _275_ sky130_fd_sc_hd__o31a_1
X_611_ _169_ _205_ _206_ vssd1 vssd1 vccd1 vccd1 _207_ sky130_fd_sc_hd__o21a_1
X_542_ net27 net10 vssd1 vssd1 vccd1 vccd1 _143_ sky130_fd_sc_hd__nand2_4
X_473_ o_csr_imm_sel o_funct3[1] o_funct3[0] _085_ vssd1 vssd1 vccd1 vccd1 o_csr_read
+ sky130_fd_sc_hd__o31a_4
X_809_ i_instruction[8] _170_ _370_ _381_ vssd1 vssd1 vccd1 vccd1 _382_ sky130_fd_sc_hd__o22a_1
X_525_ _124_ _125_ _127_ vssd1 vssd1 vccd1 vccd1 _128_ sky130_fd_sc_hd__and3_2
X_456_ o_csr_imm_sel _094_ _102_ vssd1 vssd1 vccd1 vccd1 o_imm_i[14] sky130_fd_sc_hd__a21o_2
X_387_ net29 vssd1 vssd1 vccd1 vccd1 _063_ sky130_fd_sc_hd__inv_2
X_508_ o_pc_next[13] i_pc_next[13] net21 vssd1 vssd1 vccd1 vccd1 _012_ sky130_fd_sc_hd__mux2_1
X_439_ o_rd[3] o_csr_idx[3] _092_ vssd1 vssd1 vccd1 vccd1 _097_ sky130_fd_sc_hd__mux2_1
X_790_ _159_ _365_ _362_ vssd1 vssd1 vccd1 vccd1 _366_ sky130_fd_sc_hd__o21a_1
X_842_ clknet_3_2__leaf_i_clk _011_ vssd1 vssd1 vccd1 vccd1 o_pc_next[12] sky130_fd_sc_hd__dfxtp_2
X_773_ _280_ _349_ _167_ vssd1 vssd1 vccd1 vccd1 _350_ sky130_fd_sc_hd__a21o_1
X_825_ o_pc[10] i_pc[10] net21 vssd1 vssd1 vccd1 vccd1 _057_ sky130_fd_sc_hd__mux2_1
X_756_ _163_ _166_ _187_ _334_ _193_ vssd1 vssd1 vccd1 vccd1 _335_ sky130_fd_sc_hd__a221o_1
X_687_ i_instruction[16] _126_ _145_ vssd1 vssd1 vccd1 vccd1 _274_ sky130_fd_sc_hd__mux2_1
X_610_ i_instruction[13] net9 _195_ vssd1 vssd1 vccd1 vccd1 _206_ sky130_fd_sc_hd__a21oi_1
X_541_ _141_ _142_ i_flush vssd1 vssd1 vccd1 vccd1 _017_ sky130_fd_sc_hd__a21oi_1
X_472_ o_alu_ctrl[3] net4 net1 vssd1 vssd1 vccd1 vccd1 o_imm_i[30] sky130_fd_sc_hd__a21o_2
X_808_ _074_ _132_ _187_ _122_ vssd1 vssd1 vccd1 vccd1 _381_ sky130_fd_sc_hd__o211a_1
X_739_ net26 _319_ vssd1 vssd1 vccd1 vccd1 _320_ sky130_fd_sc_hd__nand2_1
X_524_ net36 i_instruction[8] vssd1 vssd1 vccd1 vccd1 _127_ sky130_fd_sc_hd__nand2_1
X_455_ o_funct3[1] _094_ _102_ vssd1 vssd1 vccd1 vccd1 o_imm_i[13] sky130_fd_sc_hd__a21o_2
X_507_ o_pc_next[12] i_pc_next[12] net22 vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__mux2_4
X_438_ net3 _096_ vssd1 vssd1 vccd1 vccd1 o_imm_i[2] sky130_fd_sc_hd__and2_2
X_841_ clknet_3_1__leaf_i_clk _010_ vssd1 vssd1 vccd1 vccd1 o_pc_next[11] sky130_fd_sc_hd__dfxtp_2
X_772_ net37 net39 _124_ _162_ vssd1 vssd1 vccd1 vccd1 _349_ sky130_fd_sc_hd__nand4_1
X_824_ o_pc[9] i_pc[9] net22 vssd1 vssd1 vccd1 vccd1 _056_ sky130_fd_sc_hd__mux2_1
X_755_ i_instruction[10] i_instruction[11] vssd1 vssd1 vccd1 vccd1 _334_ sky130_fd_sc_hd__nand2_1
X_686_ net6 _270_ _272_ net10 vssd1 vssd1 vccd1 vccd1 _273_ sky130_fd_sc_hd__o211a_1
Xfanout1 _101_ vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_12
X_540_ net29 instruction\[1\] vssd1 vssd1 vccd1 vccd1 _142_ sky130_fd_sc_hd__nand2_1
X_471_ o_csr_idx[9] net4 net1 vssd1 vssd1 vccd1 vccd1 o_imm_i[29] sky130_fd_sc_hd__a21o_2
X_807_ net26 o_csr_idx[9] net23 _380_ vssd1 vssd1 vccd1 vccd1 _045_ sky130_fd_sc_hd__o211a_1
X_738_ net12 _316_ _318_ vssd1 vssd1 vccd1 vccd1 _319_ sky130_fd_sc_hd__o21ai_1
X_669_ i_instruction[12] _169_ vssd1 vssd1 vccd1 vccd1 _257_ sky130_fd_sc_hd__and2_2
X_523_ net36 i_instruction[8] vssd1 vssd1 vccd1 vccd1 _126_ sky130_fd_sc_hd__and2_2
X_454_ o_funct3[0] _094_ _102_ vssd1 vssd1 vccd1 vccd1 o_imm_i[12] sky130_fd_sc_hd__a21o_2
X_506_ o_pc_next[11] i_pc_next[11] net20 vssd1 vssd1 vccd1 vccd1 _010_ sky130_fd_sc_hd__mux2_1
X_437_ o_rd[2] o_csr_idx[2] _092_ vssd1 vssd1 vccd1 vccd1 _096_ sky130_fd_sc_hd__mux2_1
X_840_ clknet_3_0__leaf_i_clk _009_ vssd1 vssd1 vccd1 vccd1 o_pc_next[10] sky130_fd_sc_hd__dfxtp_2
X_771_ _340_ _347_ _165_ vssd1 vssd1 vccd1 vccd1 _348_ sky130_fd_sc_hd__o21ai_1
X_823_ o_pc[8] i_pc[8] net20 vssd1 vssd1 vccd1 vccd1 _055_ sky130_fd_sc_hd__mux2_1
X_754_ net12 _332_ _331_ net30 vssd1 vssd1 vccd1 vccd1 _333_ sky130_fd_sc_hd__a211o_1
X_685_ net5 _257_ _271_ vssd1 vssd1 vccd1 vccd1 _272_ sky130_fd_sc_hd__or3_1
Xclkbuf_3_3__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout2 net3 vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_12
X_470_ o_csr_idx[8] net4 net1 vssd1 vssd1 vccd1 vccd1 o_imm_i[28] sky130_fd_sc_hd__a21o_2
X_806_ _135_ _378_ _379_ net12 net30 vssd1 vssd1 vccd1 vccd1 _380_ sky130_fd_sc_hd__a221o_2
X_737_ _075_ _131_ _317_ net18 net11 vssd1 vssd1 vccd1 vccd1 _318_ sky130_fd_sc_hd__a221o_1
X_668_ i_flush _256_ vssd1 vssd1 vccd1 vccd1 _030_ sky130_fd_sc_hd__nor2_1
X_599_ net6 _191_ _192_ _196_ vssd1 vssd1 vccd1 vccd1 _197_ sky130_fd_sc_hd__and4_1
X_522_ net36 i_instruction[7] vssd1 vssd1 vccd1 vccd1 _125_ sky130_fd_sc_hd__nand2_2
X_453_ _079_ _101_ vssd1 vssd1 vccd1 vccd1 _102_ sky130_fd_sc_hd__and2b_4
X_505_ o_pc_next[10] i_pc_next[10] net20 vssd1 vssd1 vccd1 vccd1 _009_ sky130_fd_sc_hd__mux2_1
X_436_ _064_ _092_ _095_ vssd1 vssd1 vccd1 vccd1 o_imm_i[1] sky130_fd_sc_hd__a21oi_4
X_419_ o_csr_idx[0] _087_ vssd1 vssd1 vccd1 vccd1 o_csr_ebreak sky130_fd_sc_hd__and2_2
X_770_ _187_ net39 net34 vssd1 vssd1 vccd1 vccd1 _347_ sky130_fd_sc_hd__and3b_1
X_899_ o_csr_idx[2] vssd1 vssd1 vccd1 vccd1 o_rs2[2] sky130_fd_sc_hd__buf_2
X_822_ o_pc[7] i_pc[7] net20 vssd1 vssd1 vccd1 vccd1 _054_ sky130_fd_sc_hd__mux2_1
X_753_ _075_ _123_ net8 i_instruction[24] vssd1 vssd1 vccd1 vccd1 _332_ sky130_fd_sc_hd__a22o_1
X_684_ _126_ _164_ _168_ _131_ _218_ vssd1 vssd1 vccd1 vccd1 _271_ sky130_fd_sc_hd__o221a_1
Xfanout3 _089_ vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_12
X_805_ _120_ _122_ net8 i_instruction[29] vssd1 vssd1 vccd1 vccd1 _379_ sky130_fd_sc_hd__a22o_1
X_736_ i_instruction[22] _118_ _148_ net41 vssd1 vssd1 vccd1 vccd1 _317_ sky130_fd_sc_hd__a22o_1
X_667_ net26 _065_ _143_ _255_ vssd1 vssd1 vccd1 vccd1 _256_ sky130_fd_sc_hd__o22a_1
X_598_ _118_ _193_ vssd1 vssd1 vccd1 vccd1 _196_ sky130_fd_sc_hd__nand2_1
X_521_ i_instruction[9] i_instruction[10] i_instruction[11] net37 vssd1 vssd1 vccd1
+ vccd1 _124_ sky130_fd_sc_hd__o31ai_4
X_452_ o_csr_idx[11] net2 vssd1 vssd1 vccd1 vccd1 _101_ sky130_fd_sc_hd__and2_4
X_719_ i_instruction[20] net8 _297_ vssd1 vssd1 vccd1 vccd1 _302_ sky130_fd_sc_hd__a21o_1
X_504_ o_pc_next[9] i_pc_next[9] net22 vssd1 vssd1 vccd1 vccd1 _008_ sky130_fd_sc_hd__mux2_2
X_435_ o_rd[1] _092_ net2 vssd1 vssd1 vccd1 vccd1 _095_ sky130_fd_sc_hd__o21ai_1
X_418_ o_csr_idx[8] _086_ vssd1 vssd1 vccd1 vccd1 _087_ sky130_fd_sc_hd__nor2_4
X_898_ o_csr_idx[1] vssd1 vssd1 vccd1 vccd1 o_rs2[1] sky130_fd_sc_hd__buf_2
X_821_ o_pc[6] i_pc[6] net22 vssd1 vssd1 vccd1 vccd1 _053_ sky130_fd_sc_hd__mux2_1
X_752_ net16 _330_ vssd1 vssd1 vccd1 vccd1 _331_ sky130_fd_sc_hd__and2_1
X_683_ i_instruction[16] _172_ _269_ net14 vssd1 vssd1 vccd1 vccd1 _270_ sky130_fd_sc_hd__a22o_1
Xfanout4 _088_ vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_12
X_804_ i_instruction[29] net16 _370_ _377_ vssd1 vssd1 vccd1 vccd1 _378_ sky130_fd_sc_hd__a22o_1
X_735_ net16 _293_ _314_ _315_ vssd1 vssd1 vccd1 vccd1 _316_ sky130_fd_sc_hd__o31a_1
X_666_ net41 _173_ _241_ _254_ vssd1 vssd1 vccd1 vccd1 _255_ sky130_fd_sc_hd__o2bb2a_2
X_597_ net19 _194_ vssd1 vssd1 vccd1 vccd1 _195_ sky130_fd_sc_hd__nor2_2
X_520_ net33 i_instruction[11] vssd1 vssd1 vccd1 vccd1 _123_ sky130_fd_sc_hd__and2_2
X_451_ _079_ _099_ _100_ net2 vssd1 vssd1 vccd1 vccd1 o_imm_i[11] sky130_fd_sc_hd__o211a_2
X_718_ net15 _165_ _300_ _172_ i_instruction[20] vssd1 vssd1 vccd1 vccd1 _301_ sky130_fd_sc_hd__a32o_1
X_649_ i_instruction[12] _170_ net7 vssd1 vssd1 vccd1 vccd1 _240_ sky130_fd_sc_hd__o21a_1
X_503_ o_pc_next[8] i_pc_next[8] net20 vssd1 vssd1 vccd1 vccd1 _007_ sky130_fd_sc_hd__mux2_1
X_434_ _094_ _093_ vssd1 vssd1 vccd1 vccd1 o_imm_i[0] sky130_fd_sc_hd__and2b_2
X_417_ o_csr_imm_sel o_funct3[1] o_funct3[0] _085_ vssd1 vssd1 vccd1 vccd1 _086_ sky130_fd_sc_hd__or4b_4
X_897_ o_csr_idx[0] vssd1 vssd1 vccd1 vccd1 o_rs2[0] sky130_fd_sc_hd__buf_2
X_820_ o_pc[5] i_pc[5] net21 vssd1 vssd1 vccd1 vccd1 _052_ sky130_fd_sc_hd__mux2_1
X_751_ i_instruction[6] _136_ _172_ i_instruction[24] vssd1 vssd1 vccd1 vccd1 _330_
+ sky130_fd_sc_hd__a22o_1
X_682_ _127_ _268_ _118_ vssd1 vssd1 vccd1 vccd1 _269_ sky130_fd_sc_hd__o21ai_1
Xfanout5 _160_ vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_8
X_803_ _073_ _169_ net16 vssd1 vssd1 vccd1 vccd1 _377_ sky130_fd_sc_hd__a21oi_1
X_734_ i_instruction[4] net15 _172_ i_instruction[22] net7 vssd1 vssd1 vccd1 vccd1
+ _315_ sky130_fd_sc_hd__a221o_1
X_665_ _149_ _168_ _170_ _253_ vssd1 vssd1 vccd1 vccd1 _254_ sky130_fd_sc_hd__o211a_1
X_596_ net40 net43 net34 vssd1 vssd1 vccd1 vccd1 _194_ sky130_fd_sc_hd__o21a_2
X_450_ o_csr_idx[0] _068_ _077_ vssd1 vssd1 vccd1 vccd1 _100_ sky130_fd_sc_hd__or3b_1
X_717_ net8 _298_ _299_ _297_ vssd1 vssd1 vccd1 vccd1 _300_ sky130_fd_sc_hd__a31o_1
X_648_ net35 net43 net8 _238_ vssd1 vssd1 vccd1 vccd1 _239_ sky130_fd_sc_hd__a22o_1
X_579_ i_flush _178_ vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__nor2_1
X_502_ o_pc_next[7] i_pc_next[7] net21 vssd1 vssd1 vccd1 vccd1 _006_ sky130_fd_sc_hd__mux2_1
X_433_ _079_ _088_ vssd1 vssd1 vccd1 vccd1 _094_ sky130_fd_sc_hd__or2_4
X_416_ _066_ _080_ _084_ vssd1 vssd1 vccd1 vccd1 _085_ sky130_fd_sc_hd__nor3_4
Xclkbuf_3_6__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_896_ o_csr_idx[11] vssd1 vssd1 vccd1 vccd1 o_imm_i[31] sky130_fd_sc_hd__buf_2
X_750_ i_instruction[11] _169_ _293_ vssd1 vssd1 vccd1 vccd1 _329_ sky130_fd_sc_hd__a21o_1
X_681_ _148_ _153_ net18 _130_ vssd1 vssd1 vccd1 vccd1 _268_ sky130_fd_sc_hd__o211a_4
X_879_ clknet_3_0__leaf_i_clk _048_ vssd1 vssd1 vccd1 vccd1 o_pc[1] sky130_fd_sc_hd__dfxtp_2
Xfanout6 net7 vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_4
X_802_ net28 o_csr_idx[8] net25 _376_ vssd1 vssd1 vccd1 vccd1 _044_ sky130_fd_sc_hd__o211a_2
X_733_ net41 _192_ _149_ vssd1 vssd1 vccd1 vccd1 _314_ sky130_fd_sc_hd__a21oi_1
X_664_ i_instruction[10] _123_ _132_ _188_ vssd1 vssd1 vccd1 vccd1 _253_ sky130_fd_sc_hd__a31o_1
X_595_ net40 net43 net33 vssd1 vssd1 vccd1 vccd1 _193_ sky130_fd_sc_hd__o21ai_4
X_716_ net17 _154_ i_instruction[2] vssd1 vssd1 vccd1 vccd1 _299_ sky130_fd_sc_hd__a21o_1
X_647_ net39 _131_ _190_ vssd1 vssd1 vccd1 vccd1 _238_ sky130_fd_sc_hd__a21o_1
X_578_ _147_ _177_ net27 _068_ vssd1 vssd1 vccd1 vccd1 _178_ sky130_fd_sc_hd__o2bb2a_1
.ends

