* NGSPICE file created from rv_alu1.ext - technology: sky130A
.subckt rv_alu1
+ i_clk i_reset_n i_flush i_stall
+ i_pc[1] i_pc[2] i_pc[3] i_pc[4] i_pc[5] i_pc[6] i_pc[7] i_pc[8] i_pc[9] i_pc[10] i_pc[11] i_pc[12] i_pc[13] i_pc[14] i_pc[15] 
+ i_pc_next[1] i_pc_next[2] i_pc_next[3] i_pc_next[4] i_pc_next[5] i_pc_next[6] i_pc_next[7] i_pc_next[8] i_pc_next[9] i_pc_next[10] i_pc_next[11] i_pc_next[12] i_pc_next[13] i_pc_next[14] i_pc_next[15] 
+ i_rd[0] i_rd[1] i_rd[2] i_rd[3] i_rd[4] 
+ i_rs1[0] i_rs1[1] i_rs1[2] i_rs1[3] i_rs1[4] 
+ i_rs2[0] i_rs2[1] i_rs2[2] i_rs2[3] i_rs2[4] 
+ i_res_src[0] i_res_src[1] i_res_src[2] 
+ i_imm_i[0] i_imm_i[1] i_imm_i[2] i_imm_i[3] i_imm_i[4] i_imm_i[5] i_imm_i[6] i_imm_i[7] i_imm_i[8] i_imm_i[9] i_imm_i[10] i_imm_i[11] i_imm_i[12] i_imm_i[13] i_imm_i[14] i_imm_i[15] i_imm_i[16] i_imm_i[17] i_imm_i[18] i_imm_i[19] i_imm_i[20] i_imm_i[21] i_imm_i[22] i_imm_i[23] i_imm_i[24] i_imm_i[25] i_imm_i[26] i_imm_i[27] i_imm_i[28] i_imm_i[29] i_imm_i[30] i_imm_i[31] 
+ i_alu_ctrl[0] i_alu_ctrl[1] i_alu_ctrl[2] i_alu_ctrl[3] i_alu_ctrl[4] 
+ i_funct3[0] i_funct3[1] i_funct3[2]
+ i_reg_write i_op1_src i_op2_src i_inst_mret i_to_trap
+ i_inst_jal i_inst_jalr i_inst_branch i_inst_store 
+ i_ret_addr[1] i_ret_addr[2] i_ret_addr[3] i_ret_addr[4] i_ret_addr[5] i_ret_addr[6] i_ret_addr[7] i_ret_addr[8] i_ret_addr[9] i_ret_addr[10] i_ret_addr[11] i_ret_addr[12] i_ret_addr[13] i_ret_addr[14] i_ret_addr[15] 
+ i_reg1_data[0] i_reg1_data[1] i_reg1_data[2] i_reg1_data[3] i_reg1_data[4] i_reg1_data[5] i_reg1_data[6] i_reg1_data[7] i_reg1_data[8] i_reg1_data[9] i_reg1_data[10] i_reg1_data[11] i_reg1_data[12] i_reg1_data[13] i_reg1_data[14] i_reg1_data[15] i_reg1_data[16] i_reg1_data[17] i_reg1_data[18] i_reg1_data[19] i_reg1_data[20] i_reg1_data[21] i_reg1_data[22] i_reg1_data[23] i_reg1_data[24] i_reg1_data[25] i_reg1_data[26] i_reg1_data[27] i_reg1_data[28] i_reg1_data[29] i_reg1_data[30] i_reg1_data[31] 
+ i_reg2_data[0] i_reg2_data[1] i_reg2_data[2] i_reg2_data[3] i_reg2_data[4] i_reg2_data[5] i_reg2_data[6] i_reg2_data[7] i_reg2_data[8] i_reg2_data[9] i_reg2_data[10] i_reg2_data[11] i_reg2_data[12] i_reg2_data[13] i_reg2_data[14] i_reg2_data[15] i_reg2_data[16] i_reg2_data[17] i_reg2_data[18] i_reg2_data[19] i_reg2_data[20] i_reg2_data[21] i_reg2_data[22] i_reg2_data[23] i_reg2_data[24] i_reg2_data[25] i_reg2_data[26] i_reg2_data[27] i_reg2_data[28] i_reg2_data[29] i_reg2_data[30] i_reg2_data[31] 
+ o_op1[0] o_op1[1] o_op1[2] o_op1[3] o_op1[4] o_op1[5] o_op1[6] o_op1[7] o_op1[8] o_op1[9] o_op1[10] o_op1[11] o_op1[12] o_op1[13] o_op1[14] o_op1[15] o_op1[16] o_op1[17] o_op1[18] o_op1[19] o_op1[20] o_op1[21] o_op1[22] o_op1[23] o_op1[24] o_op1[25] o_op1[26] o_op1[27] o_op1[28] o_op1[29] o_op1[30] o_op1[31] 
+ o_op2[0] o_op2[1] o_op2[2] o_op2[3] o_op2[4] o_op2[5] o_op2[6] o_op2[7] o_op2[8] o_op2[9] o_op2[10] o_op2[11] o_op2[12] o_op2[13] o_op2[14] o_op2[15] o_op2[16] o_op2[17] o_op2[18] o_op2[19] o_op2[20] o_op2[21] o_op2[22] o_op2[23] o_op2[24] o_op2[25] o_op2[26] o_op2[27] o_op2[28] o_op2[29] o_op2[30] o_op2[31] 
+ o_store o_reg_write o_inst_jal_jalr o_inst_branch o_to_trap
+ o_alu_ctrl[0] o_alu_ctrl[1] o_alu_ctrl[2] o_alu_ctrl[3] o_alu_ctrl[4] 
+ o_rs1[0] o_rs1[1] o_rs1[2] o_rs1[3] o_rs1[4] 
+ o_rs2[0] o_rs2[1] o_rs2[2] o_rs2[3] o_rs2[4] 
+ o_rd[0] o_rd[1] o_rd[2] o_rd[3] o_rd[4] 
+ o_pc[1] o_pc[2] o_pc[3] o_pc[4] o_pc[5] o_pc[6] o_pc[7] o_pc[8] o_pc[9] o_pc[10] o_pc[11] o_pc[12] o_pc[13] o_pc[14] o_pc[15] 
+ o_pc_next[1] o_pc_next[2] o_pc_next[3] o_pc_next[4] o_pc_next[5] o_pc_next[6] o_pc_next[7] o_pc_next[8] o_pc_next[9] o_pc_next[10] o_pc_next[11] o_pc_next[12] o_pc_next[13] o_pc_next[14] o_pc_next[15] 
+ o_pc_target[1] o_pc_target[2] o_pc_target[3] o_pc_target[4] o_pc_target[5] o_pc_target[6] o_pc_target[7] o_pc_target[8] o_pc_target[9] o_pc_target[10] o_pc_target[11] o_pc_target[12] o_pc_target[13] o_pc_target[14] o_pc_target[15] 
+ o_res_src[0] o_res_src[1] o_res_src[2] 
+ o_funct3[0] o_funct3[1] o_funct3[2] 
+ vccd1 vssd1
X_432_ _109_ vssd1 vssd1 vccd1 vccd1 o_op1[9] sky130_fd_sc_hd__buf_2
X_501_ i_reg2_data[11] imm_i\[11\] _142_ vssd1 vssd1 vccd1 vccd1 _145_ sky130_fd_sc_hd__mux2_1
X_981_ clknet_3_7__leaf_i_clk _040_ vssd1 vssd1 vccd1 vccd1 o_to_trap sky130_fd_sc_hd__dfxtp_2
X_415_ _100_ vssd1 vssd1 vccd1 vccd1 o_op1[1] sky130_fd_sc_hd__buf_2
X_964_ clknet_3_5__leaf_i_clk _023_ vssd1 vssd1 vccd1 vccd1 o_funct3[1] sky130_fd_sc_hd__dfxtp_2
X_895_ _407_ vssd1 vssd1 vccd1 vccd1 _053_ sky130_fd_sc_hd__clkbuf_1
X_680_ i_rs1[2] o_rs1[2] _282_ vssd1 vssd1 vccd1 vccd1 _285_ sky130_fd_sc_hd__mux2_1
X_878_ i_pc_next[5] o_pc_next[5] _390_ vssd1 vssd1 vccd1 vccd1 _399_ sky130_fd_sc_hd__mux2_1
X_947_ clknet_3_0__leaf_i_clk _006_ vssd1 vssd1 vccd1 vccd1 op1_sel sky130_fd_sc_hd__dfxtp_2
X_801_ _288_ vssd1 vssd1 vccd1 vccd1 _354_ sky130_fd_sc_hd__clkbuf_2
X_732_ _315_ vssd1 vssd1 vccd1 vccd1 _079_ sky130_fd_sc_hd__clkbuf_1
X_663_ imm_i\[15\] _271_ vssd1 vssd1 vccd1 vccd1 _272_ sky130_fd_sc_hd__or2_1
X_594_ _174_ _208_ _210_ vssd1 vssd1 vccd1 vccd1 _211_ sky130_fd_sc_hd__a21oi_1
X_715_ i_imm_i[0] imm_i\[0\] _306_ vssd1 vssd1 vccd1 vccd1 _307_ sky130_fd_sc_hd__mux2_1
X_646_ o_pc[13] i_reg1_data[13] _168_ vssd1 vssd1 vccd1 vccd1 _257_ sky130_fd_sc_hd__mux2_1
X_577_ o_pc[5] i_reg1_data[5] inst_jalr vssd1 vssd1 vccd1 vccd1 _196_ sky130_fd_sc_hd__mux2_1
X_500_ _144_ vssd1 vssd1 vccd1 vccd1 o_op2[10] sky130_fd_sc_hd__buf_2
X_431_ i_reg1_data[9] o_pc[9] _102_ vssd1 vssd1 vccd1 vccd1 _109_ sky130_fd_sc_hd__mux2_1
X_629_ _225_ imm_i\[11\] _241_ vssd1 vssd1 vccd1 vccd1 _242_ sky130_fd_sc_hd__and3_1
X_980_ clknet_3_3__leaf_i_clk _039_ vssd1 vssd1 vccd1 vccd1 o_pc[15] sky130_fd_sc_hd__dfxtp_2
X_414_ i_reg1_data[1] o_pc[1] _099_ vssd1 vssd1 vccd1 vccd1 _100_ sky130_fd_sc_hd__mux2_1
X_963_ clknet_3_5__leaf_i_clk _022_ vssd1 vssd1 vccd1 vccd1 o_funct3[0] sky130_fd_sc_hd__dfxtp_2
X_894_ i_pc_next[13] o_pc_next[13] _281_ vssd1 vssd1 vccd1 vccd1 _407_ sky130_fd_sc_hd__mux2_1
X_946_ clknet_3_4__leaf_i_clk _005_ vssd1 vssd1 vccd1 vccd1 imm_i\[31\] sky130_fd_sc_hd__dfxtp_1
X_877_ _398_ vssd1 vssd1 vccd1 vccd1 _044_ sky130_fd_sc_hd__clkbuf_1
X_800_ _353_ vssd1 vssd1 vccd1 vccd1 _012_ sky130_fd_sc_hd__clkbuf_1
X_731_ i_imm_i[8] imm_i\[8\] _306_ vssd1 vssd1 vccd1 vccd1 _315_ sky130_fd_sc_hd__mux2_1
X_662_ o_pc[15] i_reg1_data[15] _168_ vssd1 vssd1 vccd1 vccd1 _271_ sky130_fd_sc_hd__mux2_2
X_593_ imm_i\[7\] i_ret_addr[7] inst_mret vssd1 vssd1 vccd1 vccd1 _210_ sky130_fd_sc_hd__mux2_1
X_929_ clknet_3_5__leaf_i_clk _085_ vssd1 vssd1 vccd1 vccd1 imm_i\[14\] sky130_fd_sc_hd__dfxtp_2
X_645_ imm_i\[13\] i_ret_addr[13] _167_ vssd1 vssd1 vccd1 vccd1 _256_ sky130_fd_sc_hd__mux2_1
X_714_ _281_ vssd1 vssd1 vccd1 vccd1 _306_ sky130_fd_sc_hd__clkbuf_4
X_576_ _180_ _185_ _191_ _194_ vssd1 vssd1 vccd1 vccd1 _195_ sky130_fd_sc_hd__o31a_2
X_430_ _108_ vssd1 vssd1 vccd1 vccd1 o_op1[8] sky130_fd_sc_hd__buf_2
X_628_ o_pc[11] i_reg1_data[11] _168_ vssd1 vssd1 vccd1 vccd1 _241_ sky130_fd_sc_hd__mux2_2
X_559_ _172_ _178_ _176_ _173_ vssd1 vssd1 vccd1 vccd1 _180_ sky130_fd_sc_hd__o2bb2a_2
X_413_ op1_sel vssd1 vssd1 vccd1 vccd1 _099_ sky130_fd_sc_hd__clkbuf_2
X_962_ clknet_3_6__leaf_i_clk _021_ vssd1 vssd1 vccd1 vccd1 o_reg_write sky130_fd_sc_hd__dfxtp_2
X_893_ _406_ vssd1 vssd1 vccd1 vccd1 _052_ sky130_fd_sc_hd__clkbuf_1
X_945_ clknet_3_5__leaf_i_clk _004_ vssd1 vssd1 vccd1 vccd1 imm_i\[30\] sky130_fd_sc_hd__dfxtp_1
X_876_ i_pc_next[4] o_pc_next[4] _390_ vssd1 vssd1 vccd1 vccd1 _398_ sky130_fd_sc_hd__mux2_1
X_661_ _268_ _270_ vssd1 vssd1 vccd1 vccd1 o_pc_target[14] sky130_fd_sc_hd__xnor2_4
X_592_ _170_ imm_i\[7\] _208_ vssd1 vssd1 vccd1 vccd1 _209_ sky130_fd_sc_hd__and3_1
X_730_ _314_ vssd1 vssd1 vccd1 vccd1 _078_ sky130_fd_sc_hd__clkbuf_1
X_928_ clknet_3_5__leaf_i_clk _084_ vssd1 vssd1 vccd1 vccd1 imm_i\[13\] sky130_fd_sc_hd__dfxtp_2
X_859_ _388_ vssd1 vssd1 vccd1 vccd1 _036_ sky130_fd_sc_hd__clkbuf_1
X_644_ imm_i\[13\] vssd1 vssd1 vccd1 vccd1 _255_ sky130_fd_sc_hd__inv_2
X_575_ _182_ _193_ _190_ vssd1 vssd1 vccd1 vccd1 _194_ sky130_fd_sc_hd__a21oi_1
X_713_ _305_ vssd1 vssd1 vccd1 vccd1 _070_ sky130_fd_sc_hd__clkbuf_1
X_627_ _237_ _240_ vssd1 vssd1 vccd1 vccd1 o_pc_target[10] sky130_fd_sc_hd__xnor2_4
X_558_ _172_ _179_ vssd1 vssd1 vccd1 vccd1 o_pc_target[2] sky130_fd_sc_hd__xnor2_4
X_489_ _138_ vssd1 vssd1 vccd1 vccd1 o_op2[5] sky130_fd_sc_hd__buf_2
X_412_ _098_ vssd1 vssd1 vccd1 vccd1 o_op1[0] sky130_fd_sc_hd__buf_2
X_961_ clknet_3_7__leaf_i_clk _020_ vssd1 vssd1 vccd1 vccd1 o_res_src[2] sky130_fd_sc_hd__dfxtp_2
X_892_ i_pc_next[12] o_pc_next[12] _281_ vssd1 vssd1 vccd1 vccd1 _406_ sky130_fd_sc_hd__mux2_1
X_944_ clknet_3_1__leaf_i_clk _003_ vssd1 vssd1 vccd1 vccd1 imm_i\[29\] sky130_fd_sc_hd__dfxtp_1
X_875_ _397_ vssd1 vssd1 vccd1 vccd1 _043_ sky130_fd_sc_hd__clkbuf_1
X_660_ _259_ _263_ _269_ vssd1 vssd1 vccd1 vccd1 _270_ sky130_fd_sc_hd__a21oi_2
X_591_ o_pc[7] i_reg1_data[7] inst_jalr vssd1 vssd1 vccd1 vccd1 _208_ sky130_fd_sc_hd__mux2_1
X_927_ clknet_3_5__leaf_i_clk _083_ vssd1 vssd1 vccd1 vccd1 imm_i\[12\] sky130_fd_sc_hd__dfxtp_1
X_858_ i_pc[12] o_pc[12] _379_ vssd1 vssd1 vccd1 vccd1 _388_ sky130_fd_sc_hd__mux2_1
X_789_ _346_ vssd1 vssd1 vccd1 vccd1 _008_ sky130_fd_sc_hd__clkbuf_1
X_712_ i_rs2[4] o_rs2[4] _282_ vssd1 vssd1 vccd1 vccd1 _305_ sky130_fd_sc_hd__mux2_1
X_643_ _253_ _254_ vssd1 vssd1 vccd1 vccd1 o_pc_target[12] sky130_fd_sc_hd__xnor2_4
X_574_ _186_ _187_ _188_ vssd1 vssd1 vccd1 vccd1 _193_ sky130_fd_sc_hd__a21o_1
X_626_ _238_ _232_ _239_ vssd1 vssd1 vccd1 vccd1 _240_ sky130_fd_sc_hd__o21ba_1
X_557_ _173_ _176_ _178_ vssd1 vssd1 vccd1 vccd1 _179_ sky130_fd_sc_hd__o21ai_2
X_488_ i_reg2_data[5] imm_i\[5\] _132_ vssd1 vssd1 vccd1 vccd1 _138_ sky130_fd_sc_hd__mux2_1
X_411_ _097_ i_reg1_data[0] vssd1 vssd1 vccd1 vccd1 _098_ sky130_fd_sc_hd__and2b_1
X_609_ imm_i\[9\] i_ret_addr[9] _167_ vssd1 vssd1 vccd1 vccd1 _224_ sky130_fd_sc_hd__mux2_1
X_960_ clknet_3_7__leaf_i_clk _019_ vssd1 vssd1 vccd1 vccd1 o_res_src[1] sky130_fd_sc_hd__dfxtp_2
X_891_ _405_ vssd1 vssd1 vccd1 vccd1 _051_ sky130_fd_sc_hd__clkbuf_1
X_943_ clknet_3_1__leaf_i_clk _002_ vssd1 vssd1 vccd1 vccd1 imm_i\[28\] sky130_fd_sc_hd__dfxtp_1
X_874_ i_pc_next[3] o_pc_next[3] _390_ vssd1 vssd1 vccd1 vccd1 _397_ sky130_fd_sc_hd__mux2_1
X_590_ _206_ _207_ vssd1 vssd1 vccd1 vccd1 o_pc_target[6] sky130_fd_sc_hd__xnor2_4
X_788_ _289_ _345_ vssd1 vssd1 vccd1 vccd1 _346_ sky130_fd_sc_hd__and2_1
X_926_ clknet_3_5__leaf_i_clk _082_ vssd1 vssd1 vccd1 vccd1 imm_i\[11\] sky130_fd_sc_hd__dfxtp_1
X_857_ _387_ vssd1 vssd1 vccd1 vccd1 _035_ sky130_fd_sc_hd__clkbuf_1
X_642_ _244_ _248_ _242_ vssd1 vssd1 vccd1 vccd1 _254_ sky130_fd_sc_hd__o21ba_1
X_711_ _304_ vssd1 vssd1 vccd1 vccd1 _069_ sky130_fd_sc_hd__clkbuf_1
X_573_ _191_ _192_ vssd1 vssd1 vccd1 vccd1 o_pc_target[4] sky130_fd_sc_hd__xor2_4
X_909_ clknet_3_6__leaf_i_clk _065_ vssd1 vssd1 vccd1 vccd1 o_rd[4] sky130_fd_sc_hd__dfxtp_2
X_625_ _223_ _227_ vssd1 vssd1 vccd1 vccd1 _239_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_556_ _170_ _175_ _177_ vssd1 vssd1 vccd1 vccd1 _178_ sky130_fd_sc_hd__a21o_1
X_487_ _137_ vssd1 vssd1 vccd1 vccd1 o_op2[4] sky130_fd_sc_hd__buf_2
X_410_ op1_sel vssd1 vssd1 vccd1 vccd1 _097_ sky130_fd_sc_hd__clkbuf_2
X_608_ imm_i\[9\] vssd1 vssd1 vccd1 vccd1 _223_ sky130_fd_sc_hd__inv_2
X_539_ _164_ vssd1 vssd1 vccd1 vccd1 o_op2[29] sky130_fd_sc_hd__buf_2
X_890_ i_pc_next[11] o_pc_next[11] _281_ vssd1 vssd1 vccd1 vccd1 _405_ sky130_fd_sc_hd__mux2_1
X_942_ clknet_3_1__leaf_i_clk _001_ vssd1 vssd1 vccd1 vccd1 imm_i\[27\] sky130_fd_sc_hd__dfxtp_1
X_873_ _396_ vssd1 vssd1 vccd1 vccd1 _042_ sky130_fd_sc_hd__clkbuf_1
X_925_ clknet_3_5__leaf_i_clk _081_ vssd1 vssd1 vccd1 vccd1 imm_i\[10\] sky130_fd_sc_hd__dfxtp_2
X_787_ i_inst_jal inst_jal _290_ vssd1 vssd1 vccd1 vccd1 _345_ sky130_fd_sc_hd__mux2_1
X_856_ i_pc[11] o_pc[11] _379_ vssd1 vssd1 vccd1 vccd1 _387_ sky130_fd_sc_hd__mux2_1
X_641_ _250_ _251_ _252_ vssd1 vssd1 vccd1 vccd1 _253_ sky130_fd_sc_hd__o21ba_2
X_572_ _180_ _185_ _182_ vssd1 vssd1 vccd1 vccd1 _192_ sky130_fd_sc_hd__o21ba_1
X_710_ i_rs2[3] o_rs2[3] _282_ vssd1 vssd1 vccd1 vccd1 _304_ sky130_fd_sc_hd__mux2_1
X_908_ clknet_3_3__leaf_i_clk _064_ vssd1 vssd1 vccd1 vccd1 o_rd[3] sky130_fd_sc_hd__dfxtp_2
X_839_ i_pc[3] o_pc[3] _339_ vssd1 vssd1 vccd1 vccd1 _378_ sky130_fd_sc_hd__mux2_1
X_624_ _228_ vssd1 vssd1 vccd1 vccd1 _238_ sky130_fd_sc_hd__inv_2
X_555_ imm_i\[2\] i_ret_addr[2] inst_mret vssd1 vssd1 vccd1 vccd1 _177_ sky130_fd_sc_hd__mux2_1
X_486_ i_reg2_data[4] imm_i\[4\] _132_ vssd1 vssd1 vccd1 vccd1 _137_ sky130_fd_sc_hd__mux2_1
X_607_ _220_ _222_ vssd1 vssd1 vccd1 vccd1 o_pc_target[8] sky130_fd_sc_hd__xnor2_4
X_538_ i_reg2_data[29] imm_i\[29\] op2_sel vssd1 vssd1 vccd1 vccd1 _164_ sky130_fd_sc_hd__mux2_1
X_469_ _099_ i_reg1_data[28] vssd1 vssd1 vccd1 vccd1 _128_ sky130_fd_sc_hd__and2b_1
Xclkbuf_3_2__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_941_ clknet_3_1__leaf_i_clk _000_ vssd1 vssd1 vccd1 vccd1 imm_i\[26\] sky130_fd_sc_hd__dfxtp_1
X_872_ i_pc_next[2] o_pc_next[2] _390_ vssd1 vssd1 vccd1 vccd1 _396_ sky130_fd_sc_hd__mux2_1
X_924_ clknet_3_4__leaf_i_clk _080_ vssd1 vssd1 vccd1 vccd1 imm_i\[9\] sky130_fd_sc_hd__dfxtp_2
X_786_ _344_ vssd1 vssd1 vccd1 vccd1 _007_ sky130_fd_sc_hd__clkbuf_1
X_855_ _386_ vssd1 vssd1 vccd1 vccd1 _034_ sky130_fd_sc_hd__clkbuf_1
X_640_ _225_ imm_i\[12\] _249_ vssd1 vssd1 vccd1 vccd1 _252_ sky130_fd_sc_hd__and3_1
X_571_ _189_ _190_ vssd1 vssd1 vccd1 vccd1 _191_ sky130_fd_sc_hd__or2_2
X_838_ _377_ vssd1 vssd1 vccd1 vccd1 _026_ sky130_fd_sc_hd__clkbuf_1
X_907_ clknet_3_3__leaf_i_clk _063_ vssd1 vssd1 vccd1 vccd1 o_rd[2] sky130_fd_sc_hd__dfxtp_2
X_769_ i_imm_i[26] imm_i\[26\] _328_ vssd1 vssd1 vccd1 vccd1 _335_ sky130_fd_sc_hd__mux2_1
X_623_ imm_i\[10\] _234_ _236_ vssd1 vssd1 vccd1 vccd1 _237_ sky130_fd_sc_hd__a21boi_4
X_554_ _174_ _175_ vssd1 vssd1 vccd1 vccd1 _176_ sky130_fd_sc_hd__nand2_1
X_485_ _136_ vssd1 vssd1 vccd1 vccd1 o_op2[3] sky130_fd_sc_hd__buf_2
X_606_ _211_ _215_ _221_ vssd1 vssd1 vccd1 vccd1 _222_ sky130_fd_sc_hd__o21a_1
X_468_ _127_ vssd1 vssd1 vccd1 vccd1 o_op1[27] sky130_fd_sc_hd__buf_2
X_537_ _163_ vssd1 vssd1 vccd1 vccd1 o_op2[28] sky130_fd_sc_hd__buf_2
X_940_ clknet_3_4__leaf_i_clk _096_ vssd1 vssd1 vccd1 vccd1 imm_i\[25\] sky130_fd_sc_hd__dfxtp_1
X_871_ _395_ vssd1 vssd1 vccd1 vccd1 _041_ sky130_fd_sc_hd__clkbuf_1
X_923_ clknet_3_4__leaf_i_clk _079_ vssd1 vssd1 vccd1 vccd1 imm_i\[8\] sky130_fd_sc_hd__dfxtp_1
X_854_ i_pc[10] o_pc[10] _379_ vssd1 vssd1 vccd1 vccd1 _386_ sky130_fd_sc_hd__mux2_1
X_785_ _289_ _343_ vssd1 vssd1 vccd1 vccd1 _344_ sky130_fd_sc_hd__and2_1
X_570_ imm_i\[4\] _186_ _187_ vssd1 vssd1 vccd1 vccd1 _190_ sky130_fd_sc_hd__and3_1
X_768_ _334_ vssd1 vssd1 vccd1 vccd1 _096_ sky130_fd_sc_hd__clkbuf_1
X_837_ i_pc[2] o_pc[2] _339_ vssd1 vssd1 vccd1 vccd1 _377_ sky130_fd_sc_hd__mux2_1
X_906_ clknet_3_3__leaf_i_clk _062_ vssd1 vssd1 vccd1 vccd1 o_rd[1] sky130_fd_sc_hd__dfxtp_2
X_699_ _289_ _297_ vssd1 vssd1 vccd1 vccd1 _298_ sky130_fd_sc_hd__and2_1
X_622_ _234_ _235_ vssd1 vssd1 vccd1 vccd1 _236_ sky130_fd_sc_hd__or2_1
X_484_ i_reg2_data[3] imm_i\[3\] _132_ vssd1 vssd1 vccd1 vccd1 _136_ sky130_fd_sc_hd__mux2_1
X_553_ o_pc[2] i_reg1_data[2] inst_jalr vssd1 vssd1 vccd1 vccd1 _175_ sky130_fd_sc_hd__mux2_1
X_605_ _209_ vssd1 vssd1 vccd1 vccd1 _221_ sky130_fd_sc_hd__inv_2
X_467_ _099_ i_reg1_data[27] vssd1 vssd1 vccd1 vccd1 _127_ sky130_fd_sc_hd__and2b_1
X_536_ i_reg2_data[28] imm_i\[28\] _153_ vssd1 vssd1 vccd1 vccd1 _163_ sky130_fd_sc_hd__mux2_1
X_519_ _154_ vssd1 vssd1 vccd1 vccd1 o_op2[19] sky130_fd_sc_hd__buf_2
X_870_ i_pc_next[1] o_pc_next[1] _390_ vssd1 vssd1 vccd1 vccd1 _395_ sky130_fd_sc_hd__mux2_1
X_784_ i_inst_jalr _168_ _290_ vssd1 vssd1 vccd1 vccd1 _343_ sky130_fd_sc_hd__mux2_1
X_922_ clknet_3_4__leaf_i_clk _078_ vssd1 vssd1 vccd1 vccd1 imm_i\[7\] sky130_fd_sc_hd__dfxtp_1
X_853_ _385_ vssd1 vssd1 vccd1 vccd1 _033_ sky130_fd_sc_hd__clkbuf_1
X_905_ clknet_3_3__leaf_i_clk _061_ vssd1 vssd1 vccd1 vccd1 o_rd[0] sky130_fd_sc_hd__dfxtp_2
X_767_ i_imm_i[25] imm_i\[25\] _328_ vssd1 vssd1 vccd1 vccd1 _334_ sky130_fd_sc_hd__mux2_1
X_836_ _376_ vssd1 vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__clkbuf_1
X_698_ i_rd[3] o_rd[3] _290_ vssd1 vssd1 vccd1 vccd1 _297_ sky130_fd_sc_hd__mux2_1
X_621_ imm_i\[10\] i_ret_addr[10] _167_ vssd1 vssd1 vccd1 vccd1 _235_ sky130_fd_sc_hd__mux2_1
X_552_ _170_ vssd1 vssd1 vccd1 vccd1 _174_ sky130_fd_sc_hd__buf_2
X_483_ _135_ vssd1 vssd1 vccd1 vccd1 o_op2[2] sky130_fd_sc_hd__buf_2
X_819_ _366_ vssd1 vssd1 vccd1 vccd1 _018_ sky130_fd_sc_hd__clkbuf_1
X_604_ _218_ _219_ vssd1 vssd1 vccd1 vccd1 _220_ sky130_fd_sc_hd__nor2_2
X_535_ _162_ vssd1 vssd1 vccd1 vccd1 o_op2[27] sky130_fd_sc_hd__buf_2
X_466_ _126_ vssd1 vssd1 vccd1 vccd1 o_op1[26] sky130_fd_sc_hd__buf_2
X_518_ i_reg2_data[19] imm_i\[19\] _153_ vssd1 vssd1 vccd1 vccd1 _154_ sky130_fd_sc_hd__mux2_1
X_449_ _097_ i_reg1_data[18] vssd1 vssd1 vccd1 vccd1 _118_ sky130_fd_sc_hd__and2b_1
X_921_ clknet_3_1__leaf_i_clk _077_ vssd1 vssd1 vccd1 vccd1 imm_i\[6\] sky130_fd_sc_hd__dfxtp_2
X_783_ _342_ vssd1 vssd1 vccd1 vccd1 _006_ sky130_fd_sc_hd__clkbuf_1
X_852_ i_pc[9] o_pc[9] _379_ vssd1 vssd1 vccd1 vccd1 _385_ sky130_fd_sc_hd__mux2_1
X_904_ clknet_3_2__leaf_i_clk _060_ vssd1 vssd1 vccd1 vccd1 o_rs1[4] sky130_fd_sc_hd__dfxtp_2
X_766_ _333_ vssd1 vssd1 vccd1 vccd1 _095_ sky130_fd_sc_hd__clkbuf_1
X_835_ i_pc[1] o_pc[1] _339_ vssd1 vssd1 vccd1 vccd1 _376_ sky130_fd_sc_hd__mux2_1
X_697_ _296_ vssd1 vssd1 vccd1 vccd1 _063_ sky130_fd_sc_hd__clkbuf_1
X_551_ imm_i\[2\] vssd1 vssd1 vccd1 vccd1 _173_ sky130_fd_sc_hd__inv_2
X_620_ _174_ _233_ vssd1 vssd1 vccd1 vccd1 _234_ sky130_fd_sc_hd__and2_1
Xclkbuf_3_5__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_482_ i_reg2_data[2] imm_i\[2\] _132_ vssd1 vssd1 vccd1 vccd1 _135_ sky130_fd_sc_hd__mux2_1
X_818_ _354_ _365_ vssd1 vssd1 vccd1 vccd1 _366_ sky130_fd_sc_hd__and2_1
X_749_ _324_ vssd1 vssd1 vccd1 vccd1 _087_ sky130_fd_sc_hd__clkbuf_1
X_603_ _170_ imm_i\[8\] _216_ vssd1 vssd1 vccd1 vccd1 _219_ sky130_fd_sc_hd__and3_1
X_465_ _099_ i_reg1_data[26] vssd1 vssd1 vccd1 vccd1 _126_ sky130_fd_sc_hd__and2b_1
X_534_ i_reg2_data[27] imm_i\[27\] _153_ vssd1 vssd1 vccd1 vccd1 _162_ sky130_fd_sc_hd__mux2_1
X_448_ _117_ vssd1 vssd1 vccd1 vccd1 o_op1[17] sky130_fd_sc_hd__buf_2
X_517_ op2_sel vssd1 vssd1 vccd1 vccd1 _153_ sky130_fd_sc_hd__clkbuf_4
X_851_ _384_ vssd1 vssd1 vccd1 vccd1 _032_ sky130_fd_sc_hd__clkbuf_1
X_920_ clknet_3_1__leaf_i_clk _076_ vssd1 vssd1 vccd1 vccd1 imm_i\[5\] sky130_fd_sc_hd__dfxtp_1
X_782_ i_op1_src _099_ _339_ vssd1 vssd1 vccd1 vccd1 _342_ sky130_fd_sc_hd__mux2_1
X_834_ _375_ vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__clkbuf_1
X_903_ clknet_3_2__leaf_i_clk _059_ vssd1 vssd1 vccd1 vccd1 o_rs1[3] sky130_fd_sc_hd__dfxtp_2
X_696_ _289_ _295_ vssd1 vssd1 vccd1 vccd1 _296_ sky130_fd_sc_hd__and2_1
X_765_ i_imm_i[24] imm_i\[24\] _328_ vssd1 vssd1 vccd1 vccd1 _333_ sky130_fd_sc_hd__mux2_1
X_550_ _170_ imm_i\[1\] _171_ vssd1 vssd1 vccd1 vccd1 _172_ sky130_fd_sc_hd__and3_2
X_481_ _134_ vssd1 vssd1 vccd1 vccd1 o_op2[1] sky130_fd_sc_hd__buf_2
X_817_ i_res_src[0] o_res_src[0] _351_ vssd1 vssd1 vccd1 vccd1 _365_ sky130_fd_sc_hd__mux2_1
X_748_ i_imm_i[16] imm_i\[16\] _317_ vssd1 vssd1 vccd1 vccd1 _324_ sky130_fd_sc_hd__mux2_1
X_679_ _284_ vssd1 vssd1 vccd1 vccd1 _057_ sky130_fd_sc_hd__clkbuf_1
X_602_ _174_ _216_ _217_ vssd1 vssd1 vccd1 vccd1 _218_ sky130_fd_sc_hd__a21oi_1
X_464_ _125_ vssd1 vssd1 vccd1 vccd1 o_op1[25] sky130_fd_sc_hd__buf_2
X_533_ _161_ vssd1 vssd1 vccd1 vccd1 o_op2[26] sky130_fd_sc_hd__buf_2
X_447_ _097_ i_reg1_data[17] vssd1 vssd1 vccd1 vccd1 _117_ sky130_fd_sc_hd__and2b_1
X_516_ _152_ vssd1 vssd1 vccd1 vccd1 o_op2[18] sky130_fd_sc_hd__buf_2
X_996_ clknet_3_6__leaf_i_clk _055_ vssd1 vssd1 vccd1 vccd1 o_pc_next[15] sky130_fd_sc_hd__dfxtp_2
X_781_ _341_ vssd1 vssd1 vccd1 vccd1 _005_ sky130_fd_sc_hd__clkbuf_1
X_850_ i_pc[8] o_pc[8] _379_ vssd1 vssd1 vccd1 vccd1 _384_ sky130_fd_sc_hd__mux2_1
X_979_ clknet_3_3__leaf_i_clk _038_ vssd1 vssd1 vccd1 vccd1 o_pc[14] sky130_fd_sc_hd__dfxtp_2
X_833_ i_funct3[2] o_funct3[2] _339_ vssd1 vssd1 vccd1 vccd1 _375_ sky130_fd_sc_hd__mux2_1
X_764_ _332_ vssd1 vssd1 vccd1 vccd1 _094_ sky130_fd_sc_hd__clkbuf_1
X_902_ clknet_3_2__leaf_i_clk _058_ vssd1 vssd1 vccd1 vccd1 o_rs1[2] sky130_fd_sc_hd__dfxtp_2
X_695_ i_rd[2] o_rd[2] _290_ vssd1 vssd1 vccd1 vccd1 _295_ sky130_fd_sc_hd__mux2_1
X_480_ i_reg2_data[1] imm_i\[1\] _132_ vssd1 vssd1 vccd1 vccd1 _134_ sky130_fd_sc_hd__mux2_1
X_816_ _364_ vssd1 vssd1 vccd1 vccd1 _017_ sky130_fd_sc_hd__clkbuf_1
X_747_ _323_ vssd1 vssd1 vccd1 vccd1 _086_ sky130_fd_sc_hd__clkbuf_1
X_678_ i_rs1[1] o_rs1[1] _282_ vssd1 vssd1 vccd1 vccd1 _284_ sky130_fd_sc_hd__mux2_1
X_601_ imm_i\[8\] i_ret_addr[8] inst_mret vssd1 vssd1 vccd1 vccd1 _217_ sky130_fd_sc_hd__mux2_1
X_463_ _099_ i_reg1_data[25] vssd1 vssd1 vccd1 vccd1 _125_ sky130_fd_sc_hd__and2b_1
X_532_ i_reg2_data[26] imm_i\[26\] _153_ vssd1 vssd1 vccd1 vccd1 _161_ sky130_fd_sc_hd__mux2_1
X_515_ i_reg2_data[18] imm_i\[18\] _142_ vssd1 vssd1 vccd1 vccd1 _152_ sky130_fd_sc_hd__mux2_1
X_446_ _116_ vssd1 vssd1 vccd1 vccd1 o_op1[16] sky130_fd_sc_hd__buf_2
X_995_ clknet_3_6__leaf_i_clk _054_ vssd1 vssd1 vccd1 vccd1 o_pc_next[14] sky130_fd_sc_hd__dfxtp_2
X_429_ i_reg1_data[8] o_pc[8] _102_ vssd1 vssd1 vccd1 vccd1 _108_ sky130_fd_sc_hd__mux2_1
X_780_ i_imm_i[31] imm_i\[31\] _339_ vssd1 vssd1 vccd1 vccd1 _341_ sky130_fd_sc_hd__mux2_1
X_978_ clknet_3_3__leaf_i_clk _037_ vssd1 vssd1 vccd1 vccd1 o_pc[13] sky130_fd_sc_hd__dfxtp_2
X_901_ clknet_3_2__leaf_i_clk _057_ vssd1 vssd1 vccd1 vccd1 o_rs1[1] sky130_fd_sc_hd__dfxtp_2
X_832_ _374_ vssd1 vssd1 vccd1 vccd1 _023_ sky130_fd_sc_hd__clkbuf_1
X_763_ i_imm_i[23] imm_i\[23\] _328_ vssd1 vssd1 vccd1 vccd1 _332_ sky130_fd_sc_hd__mux2_1
X_694_ _294_ vssd1 vssd1 vccd1 vccd1 _062_ sky130_fd_sc_hd__clkbuf_1
X_815_ _354_ _363_ vssd1 vssd1 vccd1 vccd1 _364_ sky130_fd_sc_hd__and2_1
X_746_ i_imm_i[15] imm_i\[15\] _317_ vssd1 vssd1 vccd1 vccd1 _323_ sky130_fd_sc_hd__mux2_1
X_677_ _283_ vssd1 vssd1 vccd1 vccd1 _056_ sky130_fd_sc_hd__clkbuf_1
X_531_ _160_ vssd1 vssd1 vccd1 vccd1 o_op2[25] sky130_fd_sc_hd__buf_2
X_600_ o_pc[8] i_reg1_data[8] inst_jalr vssd1 vssd1 vccd1 vccd1 _216_ sky130_fd_sc_hd__mux2_1
X_462_ _124_ vssd1 vssd1 vccd1 vccd1 o_op1[24] sky130_fd_sc_hd__buf_2
X_729_ i_imm_i[7] imm_i\[7\] _306_ vssd1 vssd1 vccd1 vccd1 _314_ sky130_fd_sc_hd__mux2_1
X_514_ _151_ vssd1 vssd1 vccd1 vccd1 o_op2[17] sky130_fd_sc_hd__buf_2
X_445_ _097_ i_reg1_data[16] vssd1 vssd1 vccd1 vccd1 _116_ sky130_fd_sc_hd__and2b_1
X_994_ clknet_3_6__leaf_i_clk _053_ vssd1 vssd1 vccd1 vccd1 o_pc_next[13] sky130_fd_sc_hd__dfxtp_2
X_428_ _107_ vssd1 vssd1 vccd1 vccd1 o_op1[7] sky130_fd_sc_hd__buf_2
X_977_ clknet_3_2__leaf_i_clk _036_ vssd1 vssd1 vccd1 vccd1 o_pc[12] sky130_fd_sc_hd__dfxtp_2
X_831_ i_funct3[1] o_funct3[1] _339_ vssd1 vssd1 vccd1 vccd1 _374_ sky130_fd_sc_hd__mux2_1
X_900_ clknet_3_2__leaf_i_clk _056_ vssd1 vssd1 vccd1 vccd1 o_rs1[0] sky130_fd_sc_hd__dfxtp_2
X_693_ _289_ _293_ vssd1 vssd1 vccd1 vccd1 _294_ sky130_fd_sc_hd__and2_1
X_762_ _331_ vssd1 vssd1 vccd1 vccd1 _093_ sky130_fd_sc_hd__clkbuf_1
X_814_ i_inst_store o_store _351_ vssd1 vssd1 vccd1 vccd1 _363_ sky130_fd_sc_hd__mux2_1
X_745_ _322_ vssd1 vssd1 vccd1 vccd1 _085_ sky130_fd_sc_hd__clkbuf_1
X_676_ i_rs1[0] o_rs1[0] _282_ vssd1 vssd1 vccd1 vccd1 _283_ sky130_fd_sc_hd__mux2_1
X_461_ _097_ i_reg1_data[24] vssd1 vssd1 vccd1 vccd1 _124_ sky130_fd_sc_hd__and2b_1
X_530_ i_reg2_data[25] imm_i\[25\] _153_ vssd1 vssd1 vccd1 vccd1 _160_ sky130_fd_sc_hd__mux2_1
X_659_ _255_ _258_ vssd1 vssd1 vccd1 vccd1 _269_ sky130_fd_sc_hd__nor2_1
X_728_ _313_ vssd1 vssd1 vccd1 vccd1 _077_ sky130_fd_sc_hd__clkbuf_1
X_444_ _115_ vssd1 vssd1 vccd1 vccd1 o_op1[15] sky130_fd_sc_hd__buf_2
X_513_ i_reg2_data[17] imm_i\[17\] _142_ vssd1 vssd1 vccd1 vccd1 _151_ sky130_fd_sc_hd__mux2_1
X_993_ clknet_3_6__leaf_i_clk _052_ vssd1 vssd1 vccd1 vccd1 o_pc_next[12] sky130_fd_sc_hd__dfxtp_2
X_427_ i_reg1_data[7] o_pc[7] _102_ vssd1 vssd1 vccd1 vccd1 _107_ sky130_fd_sc_hd__mux2_1
X_976_ clknet_3_2__leaf_i_clk _035_ vssd1 vssd1 vccd1 vccd1 o_pc[11] sky130_fd_sc_hd__dfxtp_2
X_830_ _373_ vssd1 vssd1 vccd1 vccd1 _022_ sky130_fd_sc_hd__clkbuf_1
X_761_ i_imm_i[22] imm_i\[22\] _328_ vssd1 vssd1 vccd1 vccd1 _331_ sky130_fd_sc_hd__mux2_1
X_692_ i_rd[1] o_rd[1] _290_ vssd1 vssd1 vccd1 vccd1 _293_ sky130_fd_sc_hd__mux2_1
X_959_ clknet_3_6__leaf_i_clk _018_ vssd1 vssd1 vccd1 vccd1 o_res_src[0] sky130_fd_sc_hd__dfxtp_2
X_813_ _362_ vssd1 vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__clkbuf_1
X_744_ i_imm_i[14] imm_i\[14\] _317_ vssd1 vssd1 vccd1 vccd1 _322_ sky130_fd_sc_hd__mux2_1
X_675_ _281_ vssd1 vssd1 vccd1 vccd1 _282_ sky130_fd_sc_hd__clkbuf_4
X_460_ _123_ vssd1 vssd1 vccd1 vccd1 o_op1[23] sky130_fd_sc_hd__buf_2
X_727_ i_imm_i[6] imm_i\[6\] _306_ vssd1 vssd1 vccd1 vccd1 _313_ sky130_fd_sc_hd__mux2_1
X_658_ _266_ _267_ vssd1 vssd1 vccd1 vccd1 _268_ sky130_fd_sc_hd__nor2_2
X_589_ _195_ _199_ _197_ vssd1 vssd1 vccd1 vccd1 _207_ sky130_fd_sc_hd__o21ba_1
X_443_ i_reg1_data[15] o_pc[15] op1_sel vssd1 vssd1 vccd1 vccd1 _115_ sky130_fd_sc_hd__mux2_1
X_512_ _150_ vssd1 vssd1 vccd1 vccd1 o_op2[16] sky130_fd_sc_hd__buf_2
X_992_ clknet_3_6__leaf_i_clk _051_ vssd1 vssd1 vccd1 vccd1 o_pc_next[11] sky130_fd_sc_hd__dfxtp_2
X_426_ _106_ vssd1 vssd1 vccd1 vccd1 o_op1[6] sky130_fd_sc_hd__buf_2
X_975_ clknet_3_2__leaf_i_clk _034_ vssd1 vssd1 vccd1 vccd1 o_pc[10] sky130_fd_sc_hd__dfxtp_2
X_760_ _330_ vssd1 vssd1 vccd1 vccd1 _092_ sky130_fd_sc_hd__clkbuf_1
X_691_ _292_ vssd1 vssd1 vccd1 vccd1 _061_ sky130_fd_sc_hd__clkbuf_1
X_958_ clknet_3_7__leaf_i_clk _017_ vssd1 vssd1 vccd1 vccd1 o_store sky130_fd_sc_hd__dfxtp_2
X_889_ _404_ vssd1 vssd1 vccd1 vccd1 _050_ sky130_fd_sc_hd__clkbuf_1
X_812_ _354_ _361_ vssd1 vssd1 vccd1 vccd1 _362_ sky130_fd_sc_hd__and2_1
X_743_ _321_ vssd1 vssd1 vccd1 vccd1 _084_ sky130_fd_sc_hd__clkbuf_1
X_674_ _280_ vssd1 vssd1 vccd1 vccd1 _281_ sky130_fd_sc_hd__clkbuf_4
X_657_ _225_ imm_i\[14\] _264_ vssd1 vssd1 vccd1 vccd1 _267_ sky130_fd_sc_hd__and3_1
X_726_ _312_ vssd1 vssd1 vccd1 vccd1 _076_ sky130_fd_sc_hd__clkbuf_1
X_588_ imm_i\[6\] _203_ _205_ vssd1 vssd1 vccd1 vccd1 _206_ sky130_fd_sc_hd__a21boi_4
X_511_ i_reg2_data[16] imm_i\[16\] _142_ vssd1 vssd1 vccd1 vccd1 _150_ sky130_fd_sc_hd__mux2_1
X_442_ _114_ vssd1 vssd1 vccd1 vccd1 o_op1[14] sky130_fd_sc_hd__buf_2
X_709_ _303_ vssd1 vssd1 vccd1 vccd1 _068_ sky130_fd_sc_hd__clkbuf_1
X_991_ clknet_3_3__leaf_i_clk _050_ vssd1 vssd1 vccd1 vccd1 o_pc_next[10] sky130_fd_sc_hd__dfxtp_2
X_425_ i_reg1_data[6] o_pc[6] _102_ vssd1 vssd1 vccd1 vccd1 _106_ sky130_fd_sc_hd__mux2_1
X_974_ clknet_3_2__leaf_i_clk _033_ vssd1 vssd1 vccd1 vccd1 o_pc[9] sky130_fd_sc_hd__dfxtp_2
X_690_ _289_ _291_ vssd1 vssd1 vccd1 vccd1 _292_ sky130_fd_sc_hd__and2_1
X_957_ clknet_3_7__leaf_i_clk _016_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[4] sky130_fd_sc_hd__dfxtp_2
X_888_ i_pc_next[10] o_pc_next[10] _281_ vssd1 vssd1 vccd1 vccd1 _404_ sky130_fd_sc_hd__mux2_1
X_811_ i_alu_ctrl[4] o_alu_ctrl[4] _351_ vssd1 vssd1 vccd1 vccd1 _361_ sky130_fd_sc_hd__mux2_1
X_742_ i_imm_i[13] imm_i\[13\] _317_ vssd1 vssd1 vccd1 vccd1 _321_ sky130_fd_sc_hd__mux2_1
X_673_ _279_ vssd1 vssd1 vccd1 vccd1 _280_ sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_3_1__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_656_ _225_ _264_ _265_ vssd1 vssd1 vccd1 vccd1 _266_ sky130_fd_sc_hd__a21oi_1
X_725_ i_imm_i[5] imm_i\[5\] _306_ vssd1 vssd1 vccd1 vccd1 _312_ sky130_fd_sc_hd__mux2_1
X_587_ _174_ _201_ _202_ _204_ vssd1 vssd1 vccd1 vccd1 _205_ sky130_fd_sc_hd__a31o_1
X_441_ i_reg1_data[14] o_pc[14] op1_sel vssd1 vssd1 vccd1 vccd1 _114_ sky130_fd_sc_hd__mux2_1
X_510_ _149_ vssd1 vssd1 vccd1 vccd1 o_op2[15] sky130_fd_sc_hd__buf_2
X_639_ imm_i\[12\] i_ret_addr[12] _167_ vssd1 vssd1 vccd1 vccd1 _251_ sky130_fd_sc_hd__mux2_1
X_708_ i_rs2[2] o_rs2[2] _282_ vssd1 vssd1 vccd1 vccd1 _303_ sky130_fd_sc_hd__mux2_1
X_990_ clknet_3_3__leaf_i_clk _049_ vssd1 vssd1 vccd1 vccd1 o_pc_next[9] sky130_fd_sc_hd__dfxtp_2
X_424_ _105_ vssd1 vssd1 vccd1 vccd1 o_op1[5] sky130_fd_sc_hd__buf_2
X_973_ clknet_3_0__leaf_i_clk _032_ vssd1 vssd1 vccd1 vccd1 o_pc[8] sky130_fd_sc_hd__dfxtp_2
X_956_ clknet_3_7__leaf_i_clk _015_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[3] sky130_fd_sc_hd__dfxtp_2
X_887_ _403_ vssd1 vssd1 vccd1 vccd1 _049_ sky130_fd_sc_hd__clkbuf_1
X_810_ _360_ vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__clkbuf_1
X_672_ i_stall i_flush i_reset_n vssd1 vssd1 vccd1 vccd1 _279_ sky130_fd_sc_hd__or3b_1
X_741_ _320_ vssd1 vssd1 vccd1 vccd1 _083_ sky130_fd_sc_hd__clkbuf_1
X_939_ clknet_3_0__leaf_i_clk _095_ vssd1 vssd1 vccd1 vccd1 imm_i\[24\] sky130_fd_sc_hd__dfxtp_1
X_724_ _311_ vssd1 vssd1 vccd1 vccd1 _075_ sky130_fd_sc_hd__clkbuf_1
X_655_ imm_i\[14\] i_ret_addr[14] _167_ vssd1 vssd1 vccd1 vccd1 _265_ sky130_fd_sc_hd__mux2_1
X_586_ imm_i\[6\] i_ret_addr[6] inst_mret vssd1 vssd1 vccd1 vccd1 _204_ sky130_fd_sc_hd__mux2_1
X_440_ _113_ vssd1 vssd1 vccd1 vccd1 o_op1[13] sky130_fd_sc_hd__buf_2
X_707_ _302_ vssd1 vssd1 vccd1 vccd1 _067_ sky130_fd_sc_hd__clkbuf_1
X_638_ _225_ _249_ vssd1 vssd1 vccd1 vccd1 _250_ sky130_fd_sc_hd__and2_1
X_569_ _186_ _187_ _188_ vssd1 vssd1 vccd1 vccd1 _189_ sky130_fd_sc_hd__a21oi_1
X_423_ i_reg1_data[5] o_pc[5] _102_ vssd1 vssd1 vccd1 vccd1 _105_ sky130_fd_sc_hd__mux2_1
X_972_ clknet_3_0__leaf_i_clk _031_ vssd1 vssd1 vccd1 vccd1 o_pc[7] sky130_fd_sc_hd__dfxtp_2
X_955_ clknet_3_7__leaf_i_clk _014_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[2] sky130_fd_sc_hd__dfxtp_2
X_886_ i_pc_next[9] o_pc_next[9] _281_ vssd1 vssd1 vccd1 vccd1 _403_ sky130_fd_sc_hd__mux2_1
X_740_ i_imm_i[12] imm_i\[12\] _317_ vssd1 vssd1 vccd1 vccd1 _320_ sky130_fd_sc_hd__mux2_1
X_671_ _172_ _278_ vssd1 vssd1 vccd1 vccd1 o_pc_target[1] sky130_fd_sc_hd__nor2_4
X_869_ _394_ vssd1 vssd1 vccd1 vccd1 _040_ sky130_fd_sc_hd__clkbuf_1
X_938_ clknet_3_0__leaf_i_clk _094_ vssd1 vssd1 vccd1 vccd1 imm_i\[23\] sky130_fd_sc_hd__dfxtp_1
X_723_ i_imm_i[4] imm_i\[4\] _306_ vssd1 vssd1 vccd1 vccd1 _311_ sky130_fd_sc_hd__mux2_1
X_654_ o_pc[14] i_reg1_data[14] _168_ vssd1 vssd1 vccd1 vccd1 _264_ sky130_fd_sc_hd__mux2_2
X_585_ _174_ _201_ _202_ vssd1 vssd1 vccd1 vccd1 _203_ sky130_fd_sc_hd__and3_1
X_637_ o_pc[12] i_reg1_data[12] _168_ vssd1 vssd1 vccd1 vccd1 _249_ sky130_fd_sc_hd__mux2_1
X_706_ i_rs2[1] o_rs2[1] _282_ vssd1 vssd1 vccd1 vccd1 _302_ sky130_fd_sc_hd__mux2_1
X_568_ imm_i\[4\] i_ret_addr[4] inst_mret vssd1 vssd1 vccd1 vccd1 _188_ sky130_fd_sc_hd__mux2_1
X_499_ i_reg2_data[10] imm_i\[10\] _142_ vssd1 vssd1 vccd1 vccd1 _144_ sky130_fd_sc_hd__mux2_1
X_422_ _104_ vssd1 vssd1 vccd1 vccd1 o_op1[4] sky130_fd_sc_hd__buf_2
X_971_ clknet_3_0__leaf_i_clk _030_ vssd1 vssd1 vccd1 vccd1 o_pc[6] sky130_fd_sc_hd__dfxtp_2
X_954_ clknet_3_7__leaf_i_clk _013_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[1] sky130_fd_sc_hd__dfxtp_2
X_885_ _402_ vssd1 vssd1 vccd1 vccd1 _048_ sky130_fd_sc_hd__clkbuf_1
X_670_ _225_ _171_ _277_ vssd1 vssd1 vccd1 vccd1 _278_ sky130_fd_sc_hd__a21oi_1
X_868_ _354_ _393_ vssd1 vssd1 vccd1 vccd1 _394_ sky130_fd_sc_hd__and2_1
X_799_ _289_ _352_ vssd1 vssd1 vccd1 vccd1 _353_ sky130_fd_sc_hd__and2_1
X_937_ clknet_3_0__leaf_i_clk _093_ vssd1 vssd1 vccd1 vccd1 imm_i\[22\] sky130_fd_sc_hd__dfxtp_1
X_653_ _259_ _263_ vssd1 vssd1 vccd1 vccd1 o_pc_target[13] sky130_fd_sc_hd__xor2_4
X_722_ _310_ vssd1 vssd1 vccd1 vccd1 _074_ sky130_fd_sc_hd__clkbuf_1
X_584_ inst_jalr o_pc[6] vssd1 vssd1 vccd1 vccd1 _202_ sky130_fd_sc_hd__or2_1
X_636_ _245_ _248_ vssd1 vssd1 vccd1 vccd1 o_pc_target[11] sky130_fd_sc_hd__xnor2_4
X_567_ inst_jalr o_pc[4] inst_mret vssd1 vssd1 vccd1 vccd1 _187_ sky130_fd_sc_hd__o21ba_1
X_705_ _301_ vssd1 vssd1 vccd1 vccd1 _066_ sky130_fd_sc_hd__clkbuf_1
X_498_ _143_ vssd1 vssd1 vccd1 vccd1 o_op2[9] sky130_fd_sc_hd__buf_2
X_421_ i_reg1_data[4] o_pc[4] _102_ vssd1 vssd1 vccd1 vccd1 _104_ sky130_fd_sc_hd__mux2_1
X_619_ o_pc[10] i_reg1_data[10] _168_ vssd1 vssd1 vccd1 vccd1 _233_ sky130_fd_sc_hd__mux2_1
X_970_ clknet_3_0__leaf_i_clk _029_ vssd1 vssd1 vccd1 vccd1 o_pc[5] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_3_4__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_953_ clknet_3_7__leaf_i_clk _012_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[0] sky130_fd_sc_hd__dfxtp_2
X_884_ i_pc_next[8] o_pc_next[8] _390_ vssd1 vssd1 vccd1 vccd1 _402_ sky130_fd_sc_hd__mux2_1
X_936_ clknet_3_0__leaf_i_clk _092_ vssd1 vssd1 vccd1 vccd1 imm_i\[21\] sky130_fd_sc_hd__dfxtp_1
X_867_ i_to_trap o_to_trap i_stall vssd1 vssd1 vccd1 vccd1 _393_ sky130_fd_sc_hd__mux2_1
X_798_ i_alu_ctrl[0] o_alu_ctrl[0] _351_ vssd1 vssd1 vccd1 vccd1 _352_ sky130_fd_sc_hd__mux2_1
X_652_ _232_ _246_ _260_ _262_ vssd1 vssd1 vccd1 vccd1 _263_ sky130_fd_sc_hd__o31ai_4
X_721_ i_imm_i[3] imm_i\[3\] _306_ vssd1 vssd1 vccd1 vccd1 _310_ sky130_fd_sc_hd__mux2_1
X_583_ i_reg1_data[6] _168_ vssd1 vssd1 vccd1 vccd1 _201_ sky130_fd_sc_hd__or2b_1
X_919_ clknet_3_1__leaf_i_clk _075_ vssd1 vssd1 vccd1 vccd1 imm_i\[4\] sky130_fd_sc_hd__dfxtp_1
X_704_ i_rs2[0] o_rs2[0] _282_ vssd1 vssd1 vccd1 vccd1 _301_ sky130_fd_sc_hd__mux2_1
X_635_ _232_ _246_ _247_ vssd1 vssd1 vccd1 vccd1 _248_ sky130_fd_sc_hd__o21ba_2
X_566_ i_reg1_data[4] inst_jalr vssd1 vssd1 vccd1 vccd1 _186_ sky130_fd_sc_hd__or2b_1
X_497_ i_reg2_data[9] imm_i\[9\] _142_ vssd1 vssd1 vccd1 vccd1 _143_ sky130_fd_sc_hd__mux2_1
X_420_ _103_ vssd1 vssd1 vccd1 vccd1 o_op1[3] sky130_fd_sc_hd__buf_2
X_618_ _228_ _232_ vssd1 vssd1 vccd1 vccd1 o_pc_target[9] sky130_fd_sc_hd__xnor2_4
X_549_ o_pc[1] i_reg1_data[1] inst_jalr vssd1 vssd1 vccd1 vccd1 _171_ sky130_fd_sc_hd__mux2_1
X_883_ _401_ vssd1 vssd1 vccd1 vccd1 _047_ sky130_fd_sc_hd__clkbuf_1
X_952_ clknet_3_0__leaf_i_clk _011_ vssd1 vssd1 vccd1 vccd1 op2_sel sky130_fd_sc_hd__dfxtp_1
X_935_ clknet_3_0__leaf_i_clk _091_ vssd1 vssd1 vccd1 vccd1 imm_i\[20\] sky130_fd_sc_hd__dfxtp_1
X_866_ _392_ vssd1 vssd1 vccd1 vccd1 _039_ sky130_fd_sc_hd__clkbuf_1
X_797_ i_stall vssd1 vssd1 vccd1 vccd1 _351_ sky130_fd_sc_hd__clkbuf_4
X_720_ _309_ vssd1 vssd1 vccd1 vccd1 _073_ sky130_fd_sc_hd__clkbuf_1
X_651_ _245_ _247_ _253_ _261_ _252_ vssd1 vssd1 vccd1 vccd1 _262_ sky130_fd_sc_hd__a311oi_4
X_582_ _195_ _200_ vssd1 vssd1 vccd1 vccd1 o_pc_target[5] sky130_fd_sc_hd__xnor2_4
X_918_ clknet_3_4__leaf_i_clk _074_ vssd1 vssd1 vccd1 vccd1 imm_i\[3\] sky130_fd_sc_hd__dfxtp_1
X_849_ _383_ vssd1 vssd1 vccd1 vccd1 _031_ sky130_fd_sc_hd__clkbuf_1
X_634_ imm_i\[10\] _234_ _236_ _239_ vssd1 vssd1 vccd1 vccd1 _247_ sky130_fd_sc_hd__a22o_1
X_703_ _300_ vssd1 vssd1 vccd1 vccd1 _065_ sky130_fd_sc_hd__clkbuf_1
X_565_ _180_ _185_ vssd1 vssd1 vccd1 vccd1 o_pc_target[3] sky130_fd_sc_hd__xor2_4
X_496_ op2_sel vssd1 vssd1 vccd1 vccd1 _142_ sky130_fd_sc_hd__clkbuf_4
X_617_ _195_ _213_ _229_ _231_ vssd1 vssd1 vccd1 vccd1 _232_ sky130_fd_sc_hd__o31a_4
X_548_ inst_mret vssd1 vssd1 vccd1 vccd1 _170_ sky130_fd_sc_hd__inv_2
X_479_ _133_ vssd1 vssd1 vccd1 vccd1 o_op2[0] sky130_fd_sc_hd__buf_2
X_951_ clknet_3_5__leaf_i_clk _010_ vssd1 vssd1 vccd1 vccd1 inst_mret sky130_fd_sc_hd__dfxtp_4
X_882_ i_pc_next[7] o_pc_next[7] _390_ vssd1 vssd1 vccd1 vccd1 _401_ sky130_fd_sc_hd__mux2_1
X_934_ clknet_3_4__leaf_i_clk _090_ vssd1 vssd1 vccd1 vccd1 imm_i\[19\] sky130_fd_sc_hd__dfxtp_1
X_796_ _350_ vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__clkbuf_1
X_865_ i_pc[15] o_pc[15] _390_ vssd1 vssd1 vccd1 vccd1 _392_ sky130_fd_sc_hd__mux2_1
X_650_ _250_ _251_ _242_ vssd1 vssd1 vccd1 vccd1 _261_ sky130_fd_sc_hd__o21a_1
X_581_ _197_ _199_ vssd1 vssd1 vccd1 vccd1 _200_ sky130_fd_sc_hd__nor2_2
X_779_ _340_ vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__clkbuf_1
X_917_ clknet_3_4__leaf_i_clk _073_ vssd1 vssd1 vccd1 vccd1 imm_i\[2\] sky130_fd_sc_hd__dfxtp_2
X_848_ i_pc[7] o_pc[7] _379_ vssd1 vssd1 vccd1 vccd1 _383_ sky130_fd_sc_hd__mux2_1
X_633_ _228_ _237_ vssd1 vssd1 vccd1 vccd1 _246_ sky130_fd_sc_hd__nand2_1
X_702_ _289_ _299_ vssd1 vssd1 vccd1 vccd1 _300_ sky130_fd_sc_hd__and2_1
X_564_ _182_ _184_ vssd1 vssd1 vccd1 vccd1 _185_ sky130_fd_sc_hd__or2_2
X_495_ _141_ vssd1 vssd1 vccd1 vccd1 o_op2[8] sky130_fd_sc_hd__buf_2
X_547_ _169_ vssd1 vssd1 vccd1 vccd1 o_inst_jal_jalr sky130_fd_sc_hd__buf_2
X_616_ _221_ _218_ _229_ _214_ _230_ vssd1 vssd1 vccd1 vccd1 _231_ sky130_fd_sc_hd__o221a_1
X_478_ i_reg2_data[0] imm_i\[0\] _132_ vssd1 vssd1 vccd1 vccd1 _133_ sky130_fd_sc_hd__mux2_1
X_950_ clknet_3_7__leaf_i_clk _009_ vssd1 vssd1 vccd1 vccd1 o_inst_branch sky130_fd_sc_hd__dfxtp_2
X_881_ _400_ vssd1 vssd1 vccd1 vccd1 _046_ sky130_fd_sc_hd__clkbuf_1
X_933_ clknet_3_4__leaf_i_clk _089_ vssd1 vssd1 vccd1 vccd1 imm_i\[18\] sky130_fd_sc_hd__dfxtp_1
X_795_ i_op2_src _132_ _339_ vssd1 vssd1 vccd1 vccd1 _350_ sky130_fd_sc_hd__mux2_1
X_864_ _391_ vssd1 vssd1 vccd1 vccd1 _038_ sky130_fd_sc_hd__clkbuf_1
X_580_ _174_ _196_ _198_ vssd1 vssd1 vccd1 vccd1 _199_ sky130_fd_sc_hd__a21oi_1
X_916_ clknet_3_1__leaf_i_clk _072_ vssd1 vssd1 vccd1 vccd1 imm_i\[1\] sky130_fd_sc_hd__dfxtp_1
X_778_ i_imm_i[30] imm_i\[30\] _339_ vssd1 vssd1 vccd1 vccd1 _340_ sky130_fd_sc_hd__mux2_1
X_847_ _382_ vssd1 vssd1 vccd1 vccd1 _030_ sky130_fd_sc_hd__clkbuf_1
X_632_ _242_ _244_ vssd1 vssd1 vccd1 vccd1 _245_ sky130_fd_sc_hd__nor2_4
X_701_ i_rd[4] o_rd[4] _290_ vssd1 vssd1 vccd1 vccd1 _299_ sky130_fd_sc_hd__mux2_1
X_563_ _174_ _181_ _183_ vssd1 vssd1 vccd1 vccd1 _184_ sky130_fd_sc_hd__a21oi_1
X_494_ i_reg2_data[8] imm_i\[8\] _132_ vssd1 vssd1 vccd1 vccd1 _141_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_7__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_546_ _167_ inst_jal _168_ vssd1 vssd1 vccd1 vccd1 _169_ sky130_fd_sc_hd__or3_1
X_615_ _219_ vssd1 vssd1 vccd1 vccd1 _230_ sky130_fd_sc_hd__inv_2
X_477_ op2_sel vssd1 vssd1 vccd1 vccd1 _132_ sky130_fd_sc_hd__clkbuf_4
X_529_ _159_ vssd1 vssd1 vccd1 vccd1 o_op2[24] sky130_fd_sc_hd__buf_2
X_880_ i_pc_next[6] o_pc_next[6] _390_ vssd1 vssd1 vccd1 vccd1 _400_ sky130_fd_sc_hd__mux2_1
X_932_ clknet_3_4__leaf_i_clk _088_ vssd1 vssd1 vccd1 vccd1 imm_i\[17\] sky130_fd_sc_hd__dfxtp_1
X_863_ i_pc[14] o_pc[14] _390_ vssd1 vssd1 vccd1 vccd1 _391_ sky130_fd_sc_hd__mux2_1
X_794_ _290_ _225_ _349_ vssd1 vssd1 vccd1 vccd1 _010_ sky130_fd_sc_hd__a21oi_1
X_915_ clknet_3_1__leaf_i_clk _071_ vssd1 vssd1 vccd1 vccd1 imm_i\[0\] sky130_fd_sc_hd__dfxtp_1
X_846_ i_pc[6] o_pc[6] _379_ vssd1 vssd1 vccd1 vccd1 _382_ sky130_fd_sc_hd__mux2_1
X_777_ _280_ vssd1 vssd1 vccd1 vccd1 _339_ sky130_fd_sc_hd__buf_4
X_700_ _298_ vssd1 vssd1 vccd1 vccd1 _064_ sky130_fd_sc_hd__clkbuf_1
X_631_ _225_ _241_ _243_ vssd1 vssd1 vccd1 vccd1 _244_ sky130_fd_sc_hd__a21oi_2
X_562_ imm_i\[3\] i_ret_addr[3] inst_mret vssd1 vssd1 vccd1 vccd1 _183_ sky130_fd_sc_hd__mux2_1
X_493_ _140_ vssd1 vssd1 vccd1 vccd1 o_op2[7] sky130_fd_sc_hd__buf_2
X_829_ i_funct3[0] o_funct3[0] _339_ vssd1 vssd1 vccd1 vccd1 _373_ sky130_fd_sc_hd__mux2_1
X_614_ _209_ _211_ _218_ _219_ vssd1 vssd1 vccd1 vccd1 _229_ sky130_fd_sc_hd__or4_1
X_476_ _131_ vssd1 vssd1 vccd1 vccd1 o_op1[31] sky130_fd_sc_hd__buf_2
X_545_ inst_jalr vssd1 vssd1 vccd1 vccd1 _168_ sky130_fd_sc_hd__buf_4
X_459_ _097_ i_reg1_data[23] vssd1 vssd1 vccd1 vccd1 _123_ sky130_fd_sc_hd__and2b_1
X_528_ i_reg2_data[24] imm_i\[24\] _153_ vssd1 vssd1 vccd1 vccd1 _159_ sky130_fd_sc_hd__mux2_1
X_931_ clknet_3_4__leaf_i_clk _087_ vssd1 vssd1 vccd1 vccd1 imm_i\[16\] sky130_fd_sc_hd__dfxtp_1
X_862_ _280_ vssd1 vssd1 vccd1 vccd1 _390_ sky130_fd_sc_hd__clkbuf_4
X_793_ _290_ i_inst_mret _289_ vssd1 vssd1 vccd1 vccd1 _349_ sky130_fd_sc_hd__o21ai_1
X_845_ _381_ vssd1 vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__clkbuf_1
X_914_ clknet_3_3__leaf_i_clk _070_ vssd1 vssd1 vccd1 vccd1 o_rs2[4] sky130_fd_sc_hd__dfxtp_2
X_776_ _338_ vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__clkbuf_1
X_630_ imm_i\[11\] i_ret_addr[11] _167_ vssd1 vssd1 vccd1 vccd1 _243_ sky130_fd_sc_hd__mux2_1
X_561_ _170_ imm_i\[3\] _181_ vssd1 vssd1 vccd1 vccd1 _182_ sky130_fd_sc_hd__and3_1
X_492_ i_reg2_data[7] imm_i\[7\] _132_ vssd1 vssd1 vccd1 vccd1 _140_ sky130_fd_sc_hd__mux2_1
X_828_ _372_ vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__clkbuf_1
X_759_ i_imm_i[21] imm_i\[21\] _328_ vssd1 vssd1 vccd1 vccd1 _330_ sky130_fd_sc_hd__mux2_1
X_613_ _223_ _224_ _227_ vssd1 vssd1 vccd1 vccd1 _228_ sky130_fd_sc_hd__mux2_2
X_544_ inst_mret vssd1 vssd1 vccd1 vccd1 _167_ sky130_fd_sc_hd__clkbuf_4
X_475_ _099_ i_reg1_data[31] vssd1 vssd1 vccd1 vccd1 _131_ sky130_fd_sc_hd__and2b_1
X_527_ _158_ vssd1 vssd1 vccd1 vccd1 o_op2[23] sky130_fd_sc_hd__buf_2
X_458_ _122_ vssd1 vssd1 vccd1 vccd1 o_op1[22] sky130_fd_sc_hd__buf_2
X_930_ clknet_3_5__leaf_i_clk _086_ vssd1 vssd1 vccd1 vccd1 imm_i\[15\] sky130_fd_sc_hd__dfxtp_2
X_792_ _348_ vssd1 vssd1 vccd1 vccd1 _009_ sky130_fd_sc_hd__clkbuf_1
X_861_ _389_ vssd1 vssd1 vccd1 vccd1 _037_ sky130_fd_sc_hd__clkbuf_1
X_913_ clknet_3_3__leaf_i_clk _069_ vssd1 vssd1 vccd1 vccd1 o_rs2[3] sky130_fd_sc_hd__dfxtp_2
X_844_ i_pc[5] o_pc[5] _379_ vssd1 vssd1 vccd1 vccd1 _381_ sky130_fd_sc_hd__mux2_1
X_775_ i_imm_i[29] imm_i\[29\] _328_ vssd1 vssd1 vccd1 vccd1 _338_ sky130_fd_sc_hd__mux2_1
X_560_ o_pc[3] i_reg1_data[3] inst_jalr vssd1 vssd1 vccd1 vccd1 _181_ sky130_fd_sc_hd__mux2_1
X_491_ _139_ vssd1 vssd1 vccd1 vccd1 o_op2[6] sky130_fd_sc_hd__buf_2
X_827_ _354_ _371_ vssd1 vssd1 vccd1 vccd1 _372_ sky130_fd_sc_hd__and2_1
X_689_ i_rd[0] o_rd[0] _290_ vssd1 vssd1 vccd1 vccd1 _291_ sky130_fd_sc_hd__mux2_1
X_758_ _329_ vssd1 vssd1 vccd1 vccd1 _091_ sky130_fd_sc_hd__clkbuf_1
X_612_ _225_ _226_ vssd1 vssd1 vccd1 vccd1 _227_ sky130_fd_sc_hd__nand2_1
X_543_ _166_ vssd1 vssd1 vccd1 vccd1 o_op2[31] sky130_fd_sc_hd__buf_2
X_474_ _130_ vssd1 vssd1 vccd1 vccd1 o_op1[30] sky130_fd_sc_hd__buf_2
X_526_ i_reg2_data[23] imm_i\[23\] _153_ vssd1 vssd1 vccd1 vccd1 _158_ sky130_fd_sc_hd__mux2_1
X_457_ _097_ i_reg1_data[22] vssd1 vssd1 vccd1 vccd1 _122_ sky130_fd_sc_hd__and2b_1
Xclkbuf_3_0__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_509_ i_reg2_data[15] imm_i\[15\] _142_ vssd1 vssd1 vccd1 vccd1 _149_ sky130_fd_sc_hd__mux2_1
X_791_ _289_ _347_ vssd1 vssd1 vccd1 vccd1 _348_ sky130_fd_sc_hd__and2_1
X_860_ i_pc[13] o_pc[13] _379_ vssd1 vssd1 vccd1 vccd1 _389_ sky130_fd_sc_hd__mux2_1
X_989_ clknet_3_6__leaf_i_clk _048_ vssd1 vssd1 vccd1 vccd1 o_pc_next[8] sky130_fd_sc_hd__dfxtp_2
X_843_ _380_ vssd1 vssd1 vccd1 vccd1 _028_ sky130_fd_sc_hd__clkbuf_1
X_912_ clknet_3_2__leaf_i_clk _068_ vssd1 vssd1 vccd1 vccd1 o_rs2[2] sky130_fd_sc_hd__dfxtp_2
X_774_ _337_ vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__clkbuf_1
X_490_ i_reg2_data[6] imm_i\[6\] _132_ vssd1 vssd1 vccd1 vccd1 _139_ sky130_fd_sc_hd__mux2_1
X_826_ i_reg_write o_reg_write _351_ vssd1 vssd1 vccd1 vccd1 _371_ sky130_fd_sc_hd__mux2_1
X_688_ i_stall vssd1 vssd1 vccd1 vccd1 _290_ sky130_fd_sc_hd__clkbuf_4
X_757_ i_imm_i[20] imm_i\[20\] _328_ vssd1 vssd1 vccd1 vccd1 _329_ sky130_fd_sc_hd__mux2_1
X_473_ _099_ i_reg1_data[30] vssd1 vssd1 vccd1 vccd1 _130_ sky130_fd_sc_hd__and2b_1
X_611_ o_pc[9] i_reg1_data[9] _168_ vssd1 vssd1 vccd1 vccd1 _226_ sky130_fd_sc_hd__mux2_1
X_542_ i_reg2_data[31] imm_i\[31\] op2_sel vssd1 vssd1 vccd1 vccd1 _166_ sky130_fd_sc_hd__mux2_1
X_809_ _354_ _359_ vssd1 vssd1 vccd1 vccd1 _360_ sky130_fd_sc_hd__and2_1
X_456_ _121_ vssd1 vssd1 vccd1 vccd1 o_op1[21] sky130_fd_sc_hd__buf_2
X_525_ _157_ vssd1 vssd1 vccd1 vccd1 o_op2[22] sky130_fd_sc_hd__buf_2
X_439_ i_reg1_data[13] o_pc[13] op1_sel vssd1 vssd1 vccd1 vccd1 _113_ sky130_fd_sc_hd__mux2_1
X_508_ _148_ vssd1 vssd1 vccd1 vccd1 o_op2[14] sky130_fd_sc_hd__buf_2
X_790_ i_inst_branch o_inst_branch _290_ vssd1 vssd1 vccd1 vccd1 _347_ sky130_fd_sc_hd__mux2_1
X_988_ clknet_3_6__leaf_i_clk _047_ vssd1 vssd1 vccd1 vccd1 o_pc_next[7] sky130_fd_sc_hd__dfxtp_2
X_842_ i_pc[4] o_pc[4] _379_ vssd1 vssd1 vccd1 vccd1 _380_ sky130_fd_sc_hd__mux2_1
X_911_ clknet_3_2__leaf_i_clk _067_ vssd1 vssd1 vccd1 vccd1 o_rs2[1] sky130_fd_sc_hd__dfxtp_2
X_773_ i_imm_i[28] imm_i\[28\] _328_ vssd1 vssd1 vccd1 vccd1 _337_ sky130_fd_sc_hd__mux2_1
X_825_ _370_ vssd1 vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__clkbuf_1
X_756_ _280_ vssd1 vssd1 vccd1 vccd1 _328_ sky130_fd_sc_hd__clkbuf_4
X_687_ _288_ vssd1 vssd1 vccd1 vccd1 _289_ sky130_fd_sc_hd__buf_2
X_610_ _174_ vssd1 vssd1 vccd1 vccd1 _225_ sky130_fd_sc_hd__buf_2
X_472_ _129_ vssd1 vssd1 vccd1 vccd1 o_op1[29] sky130_fd_sc_hd__buf_2
X_541_ _165_ vssd1 vssd1 vccd1 vccd1 o_op2[30] sky130_fd_sc_hd__buf_2
X_808_ i_alu_ctrl[3] o_alu_ctrl[3] _351_ vssd1 vssd1 vccd1 vccd1 _359_ sky130_fd_sc_hd__mux2_1
X_739_ _319_ vssd1 vssd1 vccd1 vccd1 _082_ sky130_fd_sc_hd__clkbuf_1
X_455_ _097_ i_reg1_data[21] vssd1 vssd1 vccd1 vccd1 _121_ sky130_fd_sc_hd__and2b_1
X_524_ i_reg2_data[22] imm_i\[22\] _153_ vssd1 vssd1 vccd1 vccd1 _157_ sky130_fd_sc_hd__mux2_1
X_438_ _112_ vssd1 vssd1 vccd1 vccd1 o_op1[12] sky130_fd_sc_hd__buf_2
X_507_ i_reg2_data[14] imm_i\[14\] _142_ vssd1 vssd1 vccd1 vccd1 _148_ sky130_fd_sc_hd__mux2_1
X_987_ clknet_3_6__leaf_i_clk _046_ vssd1 vssd1 vccd1 vccd1 o_pc_next[6] sky130_fd_sc_hd__dfxtp_2
X_910_ clknet_3_2__leaf_i_clk _066_ vssd1 vssd1 vccd1 vccd1 o_rs2[0] sky130_fd_sc_hd__dfxtp_2
X_841_ _280_ vssd1 vssd1 vccd1 vccd1 _379_ sky130_fd_sc_hd__clkbuf_4
X_772_ _336_ vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__clkbuf_1
X_824_ _354_ _369_ vssd1 vssd1 vccd1 vccd1 _370_ sky130_fd_sc_hd__and2_1
X_755_ _327_ vssd1 vssd1 vccd1 vccd1 _090_ sky130_fd_sc_hd__clkbuf_1
X_686_ i_flush i_reset_n vssd1 vssd1 vccd1 vccd1 _288_ sky130_fd_sc_hd__and2b_1
X_540_ i_reg2_data[30] imm_i\[30\] op2_sel vssd1 vssd1 vccd1 vccd1 _165_ sky130_fd_sc_hd__mux2_1
X_471_ _099_ i_reg1_data[29] vssd1 vssd1 vccd1 vccd1 _129_ sky130_fd_sc_hd__and2b_1
X_807_ _358_ vssd1 vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__clkbuf_1
X_669_ imm_i\[1\] i_ret_addr[1] _167_ vssd1 vssd1 vccd1 vccd1 _277_ sky130_fd_sc_hd__mux2_1
X_738_ i_imm_i[11] imm_i\[11\] _317_ vssd1 vssd1 vccd1 vccd1 _319_ sky130_fd_sc_hd__mux2_1
X_523_ _156_ vssd1 vssd1 vccd1 vccd1 o_op2[21] sky130_fd_sc_hd__buf_2
X_454_ _120_ vssd1 vssd1 vccd1 vccd1 o_op1[20] sky130_fd_sc_hd__buf_2
X_506_ _147_ vssd1 vssd1 vccd1 vccd1 o_op2[13] sky130_fd_sc_hd__buf_2
X_437_ i_reg1_data[12] o_pc[12] _102_ vssd1 vssd1 vccd1 vccd1 _112_ sky130_fd_sc_hd__mux2_1
X_986_ clknet_3_6__leaf_i_clk _045_ vssd1 vssd1 vccd1 vccd1 o_pc_next[5] sky130_fd_sc_hd__dfxtp_2
X_840_ _378_ vssd1 vssd1 vccd1 vccd1 _027_ sky130_fd_sc_hd__clkbuf_1
X_771_ i_imm_i[27] imm_i\[27\] _328_ vssd1 vssd1 vccd1 vccd1 _336_ sky130_fd_sc_hd__mux2_1
X_969_ clknet_3_0__leaf_i_clk _028_ vssd1 vssd1 vccd1 vccd1 o_pc[4] sky130_fd_sc_hd__dfxtp_4
X_823_ i_res_src[2] o_res_src[2] _351_ vssd1 vssd1 vccd1 vccd1 _369_ sky130_fd_sc_hd__mux2_1
X_754_ i_imm_i[19] imm_i\[19\] _317_ vssd1 vssd1 vccd1 vccd1 _327_ sky130_fd_sc_hd__mux2_1
X_685_ _287_ vssd1 vssd1 vccd1 vccd1 _060_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_3__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_470_ _128_ vssd1 vssd1 vccd1 vccd1 o_op1[28] sky130_fd_sc_hd__buf_2
X_806_ _354_ _357_ vssd1 vssd1 vccd1 vccd1 _358_ sky130_fd_sc_hd__and2_1
X_668_ _274_ _276_ vssd1 vssd1 vccd1 vccd1 o_pc_target[15] sky130_fd_sc_hd__xnor2_4
X_737_ _318_ vssd1 vssd1 vccd1 vccd1 _081_ sky130_fd_sc_hd__clkbuf_1
X_599_ _212_ _215_ vssd1 vssd1 vccd1 vccd1 o_pc_target[7] sky130_fd_sc_hd__xnor2_4
X_453_ _097_ i_reg1_data[20] vssd1 vssd1 vccd1 vccd1 _120_ sky130_fd_sc_hd__and2b_1
X_522_ i_reg2_data[21] imm_i\[21\] _153_ vssd1 vssd1 vccd1 vccd1 _156_ sky130_fd_sc_hd__mux2_1
X_436_ _111_ vssd1 vssd1 vccd1 vccd1 o_op1[11] sky130_fd_sc_hd__buf_2
X_505_ i_reg2_data[13] imm_i\[13\] _142_ vssd1 vssd1 vccd1 vccd1 _147_ sky130_fd_sc_hd__mux2_1
X_985_ clknet_3_3__leaf_i_clk _044_ vssd1 vssd1 vccd1 vccd1 o_pc_next[4] sky130_fd_sc_hd__dfxtp_2
X_419_ i_reg1_data[3] o_pc[3] _102_ vssd1 vssd1 vccd1 vccd1 _103_ sky130_fd_sc_hd__mux2_1
X_770_ _335_ vssd1 vssd1 vccd1 vccd1 _000_ sky130_fd_sc_hd__clkbuf_1
X_968_ clknet_3_0__leaf_i_clk _027_ vssd1 vssd1 vccd1 vccd1 o_pc[3] sky130_fd_sc_hd__dfxtp_2
X_899_ _409_ vssd1 vssd1 vccd1 vccd1 _055_ sky130_fd_sc_hd__clkbuf_1
X_822_ _368_ vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__clkbuf_1
X_753_ _326_ vssd1 vssd1 vccd1 vccd1 _089_ sky130_fd_sc_hd__clkbuf_1
X_684_ i_rs1[4] o_rs1[4] _282_ vssd1 vssd1 vccd1 vccd1 _287_ sky130_fd_sc_hd__mux2_1
X_805_ i_alu_ctrl[2] o_alu_ctrl[2] _351_ vssd1 vssd1 vccd1 vccd1 _357_ sky130_fd_sc_hd__mux2_1
X_736_ i_imm_i[10] imm_i\[10\] _317_ vssd1 vssd1 vccd1 vccd1 _318_ sky130_fd_sc_hd__mux2_1
X_667_ _266_ _275_ vssd1 vssd1 vccd1 vccd1 _276_ sky130_fd_sc_hd__or2_2
X_598_ _195_ _213_ _214_ vssd1 vssd1 vccd1 vccd1 _215_ sky130_fd_sc_hd__o21a_1
X_452_ _119_ vssd1 vssd1 vccd1 vccd1 o_op1[19] sky130_fd_sc_hd__buf_2
X_521_ _155_ vssd1 vssd1 vccd1 vccd1 o_op2[20] sky130_fd_sc_hd__buf_2
X_719_ i_imm_i[2] imm_i\[2\] _306_ vssd1 vssd1 vccd1 vccd1 _309_ sky130_fd_sc_hd__mux2_1
X_435_ i_reg1_data[11] o_pc[11] _102_ vssd1 vssd1 vccd1 vccd1 _111_ sky130_fd_sc_hd__mux2_1
X_504_ _146_ vssd1 vssd1 vccd1 vccd1 o_op2[12] sky130_fd_sc_hd__buf_2
X_984_ clknet_3_3__leaf_i_clk _043_ vssd1 vssd1 vccd1 vccd1 o_pc_next[3] sky130_fd_sc_hd__dfxtp_2
X_418_ op1_sel vssd1 vssd1 vccd1 vccd1 _102_ sky130_fd_sc_hd__clkbuf_4
X_898_ i_pc_next[15] o_pc_next[15] _281_ vssd1 vssd1 vccd1 vccd1 _409_ sky130_fd_sc_hd__mux2_1
X_967_ clknet_3_1__leaf_i_clk _026_ vssd1 vssd1 vccd1 vccd1 o_pc[2] sky130_fd_sc_hd__dfxtp_2
X_821_ _354_ _367_ vssd1 vssd1 vccd1 vccd1 _368_ sky130_fd_sc_hd__and2_1
X_752_ i_imm_i[18] imm_i\[18\] _317_ vssd1 vssd1 vccd1 vccd1 _326_ sky130_fd_sc_hd__mux2_1
X_683_ _286_ vssd1 vssd1 vccd1 vccd1 _059_ sky130_fd_sc_hd__clkbuf_1
X_804_ _356_ vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__clkbuf_1
X_735_ _281_ vssd1 vssd1 vccd1 vccd1 _317_ sky130_fd_sc_hd__clkbuf_4
X_666_ _259_ _263_ _267_ _269_ vssd1 vssd1 vccd1 vccd1 _275_ sky130_fd_sc_hd__a211oi_1
X_597_ imm_i\[6\] _203_ _205_ _197_ vssd1 vssd1 vccd1 vccd1 _214_ sky130_fd_sc_hd__a22oi_2
X_520_ i_reg2_data[20] imm_i\[20\] _153_ vssd1 vssd1 vccd1 vccd1 _155_ sky130_fd_sc_hd__mux2_1
X_451_ _097_ i_reg1_data[19] vssd1 vssd1 vccd1 vccd1 _119_ sky130_fd_sc_hd__and2b_1
X_649_ _245_ _253_ vssd1 vssd1 vccd1 vccd1 _260_ sky130_fd_sc_hd__nand2_1
X_718_ _308_ vssd1 vssd1 vccd1 vccd1 _072_ sky130_fd_sc_hd__clkbuf_1
X_503_ i_reg2_data[12] imm_i\[12\] _142_ vssd1 vssd1 vccd1 vccd1 _146_ sky130_fd_sc_hd__mux2_1
X_434_ _110_ vssd1 vssd1 vccd1 vccd1 o_op1[10] sky130_fd_sc_hd__buf_2
X_983_ clknet_3_3__leaf_i_clk _042_ vssd1 vssd1 vccd1 vccd1 o_pc_next[2] sky130_fd_sc_hd__dfxtp_2
X_417_ _101_ vssd1 vssd1 vccd1 vccd1 o_op1[2] sky130_fd_sc_hd__buf_2
X_897_ _408_ vssd1 vssd1 vccd1 vccd1 _054_ sky130_fd_sc_hd__clkbuf_1
X_966_ clknet_3_1__leaf_i_clk _025_ vssd1 vssd1 vccd1 vccd1 o_pc[1] sky130_fd_sc_hd__dfxtp_2
X_820_ i_res_src[1] o_res_src[1] _351_ vssd1 vssd1 vccd1 vccd1 _367_ sky130_fd_sc_hd__mux2_1
X_751_ _325_ vssd1 vssd1 vccd1 vccd1 _088_ sky130_fd_sc_hd__clkbuf_1
X_682_ i_rs1[3] o_rs1[3] _282_ vssd1 vssd1 vccd1 vccd1 _286_ sky130_fd_sc_hd__mux2_1
X_949_ clknet_3_5__leaf_i_clk _008_ vssd1 vssd1 vccd1 vccd1 inst_jal sky130_fd_sc_hd__dfxtp_1
X_803_ _354_ _355_ vssd1 vssd1 vccd1 vccd1 _356_ sky130_fd_sc_hd__and2_1
X_665_ _167_ i_ret_addr[15] _272_ _273_ vssd1 vssd1 vccd1 vccd1 _274_ sky130_fd_sc_hd__a22o_2
X_734_ _316_ vssd1 vssd1 vccd1 vccd1 _080_ sky130_fd_sc_hd__clkbuf_1
X_596_ _200_ _206_ vssd1 vssd1 vccd1 vccd1 _213_ sky130_fd_sc_hd__nand2_1
X_450_ _118_ vssd1 vssd1 vccd1 vccd1 o_op1[18] sky130_fd_sc_hd__buf_2
X_648_ _255_ _256_ _258_ vssd1 vssd1 vccd1 vccd1 _259_ sky130_fd_sc_hd__mux2_2
X_717_ i_imm_i[1] imm_i\[1\] _306_ vssd1 vssd1 vccd1 vccd1 _308_ sky130_fd_sc_hd__mux2_1
X_579_ imm_i\[5\] i_ret_addr[5] inst_mret vssd1 vssd1 vccd1 vccd1 _198_ sky130_fd_sc_hd__mux2_1
X_433_ i_reg1_data[10] o_pc[10] _102_ vssd1 vssd1 vccd1 vccd1 _110_ sky130_fd_sc_hd__mux2_1
X_502_ _145_ vssd1 vssd1 vccd1 vccd1 o_op2[11] sky130_fd_sc_hd__buf_2
X_982_ clknet_3_3__leaf_i_clk _041_ vssd1 vssd1 vccd1 vccd1 o_pc_next[1] sky130_fd_sc_hd__dfxtp_2
X_416_ i_reg1_data[2] o_pc[2] _099_ vssd1 vssd1 vccd1 vccd1 _101_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6__f_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_965_ clknet_3_5__leaf_i_clk _024_ vssd1 vssd1 vccd1 vccd1 o_funct3[2] sky130_fd_sc_hd__dfxtp_2
X_896_ i_pc_next[14] o_pc_next[14] _281_ vssd1 vssd1 vccd1 vccd1 _408_ sky130_fd_sc_hd__mux2_1
X_750_ i_imm_i[17] imm_i\[17\] _317_ vssd1 vssd1 vccd1 vccd1 _325_ sky130_fd_sc_hd__mux2_1
X_681_ _285_ vssd1 vssd1 vccd1 vccd1 _058_ sky130_fd_sc_hd__clkbuf_1
X_948_ clknet_3_5__leaf_i_clk _007_ vssd1 vssd1 vccd1 vccd1 inst_jalr sky130_fd_sc_hd__dfxtp_4
X_879_ _399_ vssd1 vssd1 vccd1 vccd1 _045_ sky130_fd_sc_hd__clkbuf_1
X_802_ i_alu_ctrl[1] o_alu_ctrl[1] _351_ vssd1 vssd1 vccd1 vccd1 _355_ sky130_fd_sc_hd__mux2_1
X_664_ imm_i\[15\] _271_ _167_ vssd1 vssd1 vccd1 vccd1 _273_ sky130_fd_sc_hd__a21oi_1
X_733_ i_imm_i[9] imm_i\[9\] _306_ vssd1 vssd1 vccd1 vccd1 _316_ sky130_fd_sc_hd__mux2_1
X_595_ _209_ _211_ vssd1 vssd1 vccd1 vccd1 _212_ sky130_fd_sc_hd__nor2_2
X_716_ _307_ vssd1 vssd1 vccd1 vccd1 _071_ sky130_fd_sc_hd__clkbuf_1
X_647_ _225_ _257_ vssd1 vssd1 vccd1 vccd1 _258_ sky130_fd_sc_hd__nand2_1
X_578_ _174_ imm_i\[5\] _196_ vssd1 vssd1 vccd1 vccd1 _197_ sky130_fd_sc_hd__and3_1
.ends
