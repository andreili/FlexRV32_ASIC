
.include ../../elements/inc_lib.spice
.include simulation/rv_fetch_buf.spice

.param VCC=1.8

VVCC VCC 0 PWL 0ns 0 1ns 0 1.1ns {VCC}
Vi_clk i_clk 0 PULSE 0 {VCC} 10ps 20ps 20ps 960ps 2000ps
VVSS VSS 0 PWL 0n 0

.include simulation/stimuli_rv_fetch_buf.cir
.options timeint reltol=1e-3 abstol=1e-5
.options linsol type=belos AZ_tol=1.0e-3
.tran 1p 4n
.print tran format=raw file=simulation/rv_fetch_buf.spice.raw v(*)

.GLOBAL VCC
.GLOBAL VSS
.end
