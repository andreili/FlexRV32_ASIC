
.include ../../elements/inc_lib.spice

.param VCC=1.8

VVCC VCC 0 PWL 0ns 0 1ns 0 1.1ns {VCC}
VVSS VSS 0 PWL 0n 0

.OPTIONS MEASURE MEASFAIL=1
.OPTIONS LINSOL type=klu2 AZ_tol=1.0e-3 TR_PARTITION=1 TR_PARTITION_TYPE=GRAPH
.OPTIONS TIMEINT RELTOL=1e-3 ABSTOL=1e-5 method=gear
.OPTIONS DIST STRATEGY=2

.GLOBAL VCC
.GLOBAL VSS
