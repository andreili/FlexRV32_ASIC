
.include ../block_head.spice
.include simulation/rom.spice

.include simulation/stimuli_rom.cir

.tran 1p 200n
.print tran format=raw file=simulation/rom.spice.raw v(*) i(*)

*.meas tran rd_v_0[*] find v(rd[*]) at=1.8n

.meas tran power avg par('(-1*v(VCC)*I(VVCC))') from=1.4n to=19n

.end
