** sch_path: /media/FlexRV32/asic/blocks/rv_decode_comp/rv_decode_comp.sch
**.subckt rv_decode_comp o_illegal_instruction
*+ o_instruction[31],o_instruction[30],o_instruction[29],o_instruction[28],o_instruction[27],o_instruction[26],o_instruction[25],o_instruction[24],o_instruction[23],o_instruction[22],o_instruction[21],o_instruction[20],o_instruction[19],o_instruction[18],o_instruction[17],o_instruction[16],o_instruction[15],o_instruction[14],o_instruction[13],o_instruction[12],o_instruction[11],o_instruction[10],o_instruction[9],o_instruction[8],o_instruction[7],o_instruction[6],o_instruction[5],o_instruction[4],o_instruction[3],o_instruction[2],o_instruction[1],o_instruction[0]
*+ i_instruction[31],i_instruction[30],i_instruction[29],i_instruction[28],i_instruction[27],i_instruction[26],i_instruction[25],i_instruction[24],i_instruction[23],i_instruction[22],i_instruction[21],i_instruction[20],i_instruction[19],i_instruction[18],i_instruction[17],i_instruction[16],i_instruction[15],i_instruction[14],i_instruction[13],i_instruction[12],i_instruction[11],i_instruction[10],i_instruction[9],i_instruction[8],i_instruction[7],i_instruction[6],i_instruction[5],i_instruction[4],i_instruction[3],i_instruction[2],i_instruction[1],i_instruction[0]
*.opin o_illegal_instruction
*.opin
*+ o_instruction[31],o_instruction[30],o_instruction[29],o_instruction[28],o_instruction[27],o_instruction[26],o_instruction[25],o_instruction[24],o_instruction[23],o_instruction[22],o_instruction[21],o_instruction[20],o_instruction[19],o_instruction[18],o_instruction[17],o_instruction[16],o_instruction[15],o_instruction[14],o_instruction[13],o_instruction[12],o_instruction[11],o_instruction[10],o_instruction[9],o_instruction[8],o_instruction[7],o_instruction[6],o_instruction[5],o_instruction[4],o_instruction[3],o_instruction[2],o_instruction[1],o_instruction[0]
*.ipin
*+ i_instruction[31],i_instruction[30],i_instruction[29],i_instruction[28],i_instruction[27],i_instruction[26],i_instruction[25],i_instruction[24],i_instruction[23],i_instruction[22],i_instruction[21],i_instruction[20],i_instruction[19],i_instruction[18],i_instruction[17],i_instruction[16],i_instruction[15],i_instruction[14],i_instruction[13],i_instruction[12],i_instruction[11],i_instruction[10],i_instruction[9],i_instruction[8],i_instruction[7],i_instruction[6],i_instruction[5],i_instruction[4],i_instruction[3],i_instruction[2],i_instruction[1],i_instruction[0]
x1[32] i_instruction[1] net4[32] o_illegal_instruction net1 net5[32] mux2
x1[31] i_instruction[1] net4[31] o_instruction[31] net1 net5[31] mux2
x1[30] i_instruction[1] net4[30] o_instruction[30] net1 net5[30] mux2
x1[29] i_instruction[1] net4[29] o_instruction[29] net1 net5[29] mux2
x1[28] i_instruction[1] net4[28] o_instruction[28] net1 net5[28] mux2
x1[27] i_instruction[1] net4[27] o_instruction[27] net1 net5[27] mux2
x1[26] i_instruction[1] net4[26] o_instruction[26] net1 net5[26] mux2
x1[25] i_instruction[1] net4[25] o_instruction[25] net1 net5[25] mux2
x1[24] i_instruction[1] net4[24] o_instruction[24] net1 net5[24] mux2
x1[23] i_instruction[1] net4[23] o_instruction[23] net1 net5[23] mux2
x1[22] i_instruction[1] net4[22] o_instruction[22] net1 net5[22] mux2
x1[21] i_instruction[1] net4[21] o_instruction[21] net1 net5[21] mux2
x1[20] i_instruction[1] net4[20] o_instruction[20] net1 net5[20] mux2
x1[19] i_instruction[1] net4[19] o_instruction[19] net1 net5[19] mux2
x1[18] i_instruction[1] net4[18] o_instruction[18] net1 net5[18] mux2
x1[17] i_instruction[1] net4[17] o_instruction[17] net1 net5[17] mux2
x1[16] i_instruction[1] net4[16] o_instruction[16] net1 net5[16] mux2
x1[15] i_instruction[1] net4[15] o_instruction[15] net1 net5[15] mux2
x1[14] i_instruction[1] net4[14] o_instruction[14] net1 net5[14] mux2
x1[13] i_instruction[1] net4[13] o_instruction[13] net1 net5[13] mux2
x1[12] i_instruction[1] net4[12] o_instruction[12] net1 net5[12] mux2
x1[11] i_instruction[1] net4[11] o_instruction[11] net1 net5[11] mux2
x1[10] i_instruction[1] net4[10] o_instruction[10] net1 net5[10] mux2
x1[9] i_instruction[1] net4[9] o_instruction[9] net1 net5[9] mux2
x1[8] i_instruction[1] net4[8] o_instruction[8] net1 net5[8] mux2
x1[7] i_instruction[1] net4[7] o_instruction[7] net1 net5[7] mux2
x1[6] i_instruction[1] net4[6] o_instruction[6] net1 net5[6] mux2
x1[5] i_instruction[1] net4[5] o_instruction[5] net1 net5[5] mux2
x1[4] i_instruction[1] net4[4] o_instruction[4] net1 net5[4] mux2
x1[3] i_instruction[1] net4[3] o_instruction[3] net1 net5[3] mux2
x1[2] i_instruction[1] net4[2] o_instruction[2] net1 net5[2] mux2
x1[1] i_instruction[1] net4[1] o_instruction[1] net1 net5[1] mux2
x1[0] i_instruction[1] net4[0] o_instruction[0] net1 net5[0] mux2
x1 i_instruction[1] VSS VSS VCC VCC net1 sky130_fd_sc_hd__inv_1
x2[32] i_instruction[0] VCC net4[32] net2 net47[32] mux2
x2[31] i_instruction[0] i_instruction[31] net4[31] net2 net47[31] mux2
x2[30] i_instruction[0] i_instruction[30] net4[30] net2 net47[30] mux2
x2[29] i_instruction[0] i_instruction[29] net4[29] net2 net47[29] mux2
x2[28] i_instruction[0] i_instruction[28] net4[28] net2 net47[28] mux2
x2[27] i_instruction[0] i_instruction[27] net4[27] net2 net47[27] mux2
x2[26] i_instruction[0] i_instruction[26] net4[26] net2 net47[26] mux2
x2[25] i_instruction[0] i_instruction[25] net4[25] net2 net47[25] mux2
x2[24] i_instruction[0] i_instruction[24] net4[24] net2 net47[24] mux2
x2[23] i_instruction[0] i_instruction[23] net4[23] net2 net47[23] mux2
x2[22] i_instruction[0] i_instruction[22] net4[22] net2 net47[22] mux2
x2[21] i_instruction[0] i_instruction[21] net4[21] net2 net47[21] mux2
x2[20] i_instruction[0] i_instruction[20] net4[20] net2 net47[20] mux2
x2[19] i_instruction[0] i_instruction[19] net4[19] net2 net47[19] mux2
x2[18] i_instruction[0] i_instruction[18] net4[18] net2 net47[18] mux2
x2[17] i_instruction[0] i_instruction[17] net4[17] net2 net47[17] mux2
x2[16] i_instruction[0] i_instruction[16] net4[16] net2 net47[16] mux2
x2[15] i_instruction[0] i_instruction[15] net4[15] net2 net47[15] mux2
x2[14] i_instruction[0] i_instruction[14] net4[14] net2 net47[14] mux2
x2[13] i_instruction[0] i_instruction[13] net4[13] net2 net47[13] mux2
x2[12] i_instruction[0] i_instruction[12] net4[12] net2 net47[12] mux2
x2[11] i_instruction[0] i_instruction[11] net4[11] net2 net47[11] mux2
x2[10] i_instruction[0] i_instruction[10] net4[10] net2 net47[10] mux2
x2[9] i_instruction[0] i_instruction[9] net4[9] net2 net47[9] mux2
x2[8] i_instruction[0] i_instruction[8] net4[8] net2 net47[8] mux2
x2[7] i_instruction[0] i_instruction[7] net4[7] net2 net47[7] mux2
x2[6] i_instruction[0] i_instruction[6] net4[6] net2 net47[6] mux2
x2[5] i_instruction[0] i_instruction[5] net4[5] net2 net47[5] mux2
x2[4] i_instruction[0] i_instruction[4] net4[4] net2 net47[4] mux2
x2[3] i_instruction[0] i_instruction[3] net4[3] net2 net47[3] mux2
x2[2] i_instruction[0] i_instruction[2] net4[2] net2 net47[2] mux2
x2[1] i_instruction[0] i_instruction[1] net4[1] net2 net47[1] mux2
x2[0] i_instruction[0] i_instruction[0] net4[0] net2 net47[0] mux2
x3 i_instruction[0] VSS VSS VCC VCC net2 sky130_fd_sc_hd__inv_1
x3[32] i_instruction[0] net18[32] net5[32] net3 net7[32] mux2
x3[31] i_instruction[0] net18[31] net5[31] net3 net7[31] mux2
x3[30] i_instruction[0] net18[30] net5[30] net3 net7[30] mux2
x3[29] i_instruction[0] net18[29] net5[29] net3 net7[29] mux2
x3[28] i_instruction[0] net18[28] net5[28] net3 net7[28] mux2
x3[27] i_instruction[0] net18[27] net5[27] net3 net7[27] mux2
x3[26] i_instruction[0] net18[26] net5[26] net3 net7[26] mux2
x3[25] i_instruction[0] net18[25] net5[25] net3 net7[25] mux2
x3[24] i_instruction[0] net18[24] net5[24] net3 net7[24] mux2
x3[23] i_instruction[0] net18[23] net5[23] net3 net7[23] mux2
x3[22] i_instruction[0] net18[22] net5[22] net3 net7[22] mux2
x3[21] i_instruction[0] net18[21] net5[21] net3 net7[21] mux2
x3[20] i_instruction[0] net18[20] net5[20] net3 net7[20] mux2
x3[19] i_instruction[0] net18[19] net5[19] net3 net7[19] mux2
x3[18] i_instruction[0] net18[18] net5[18] net3 net7[18] mux2
x3[17] i_instruction[0] net18[17] net5[17] net3 net7[17] mux2
x3[16] i_instruction[0] net18[16] net5[16] net3 net7[16] mux2
x3[15] i_instruction[0] net18[15] net5[15] net3 net7[15] mux2
x3[14] i_instruction[0] net18[14] net5[14] net3 net7[14] mux2
x3[13] i_instruction[0] net18[13] net5[13] net3 net7[13] mux2
x3[12] i_instruction[0] net18[12] net5[12] net3 net7[12] mux2
x3[11] i_instruction[0] net18[11] net5[11] net3 net7[11] mux2
x3[10] i_instruction[0] net18[10] net5[10] net3 net7[10] mux2
x3[9] i_instruction[0] net18[9] net5[9] net3 net7[9] mux2
x3[8] i_instruction[0] net18[8] net5[8] net3 net7[8] mux2
x3[7] i_instruction[0] net18[7] net5[7] net3 net7[7] mux2
x3[6] i_instruction[0] net18[6] net5[6] net3 net7[6] mux2
x3[5] i_instruction[0] net18[5] net5[5] net3 net7[5] mux2
x3[4] i_instruction[0] net18[4] net5[4] net3 net7[4] mux2
x3[3] i_instruction[0] net18[3] net5[3] net3 net7[3] mux2
x3[2] i_instruction[0] net18[2] net5[2] net3 net7[2] mux2
x3[1] i_instruction[0] net18[1] net5[1] net3 net7[1] mux2
x3[0] i_instruction[0] net18[0] net5[0] net3 net7[0] mux2
x4 i_instruction[0] VSS VSS VCC VCC net3 sky130_fd_sc_hd__inv_1
x4[32] i_instruction[15] net11[32] net7[32] net6 net9[32] mux2
x4[31] i_instruction[15] net11[31] net7[31] net6 net9[31] mux2
x4[30] i_instruction[15] net11[30] net7[30] net6 net9[30] mux2
x4[29] i_instruction[15] net11[29] net7[29] net6 net9[29] mux2
x4[28] i_instruction[15] net11[28] net7[28] net6 net9[28] mux2
x4[27] i_instruction[15] net11[27] net7[27] net6 net9[27] mux2
x4[26] i_instruction[15] net11[26] net7[26] net6 net9[26] mux2
x4[25] i_instruction[15] net11[25] net7[25] net6 net9[25] mux2
x4[24] i_instruction[15] net11[24] net7[24] net6 net9[24] mux2
x4[23] i_instruction[15] net11[23] net7[23] net6 net9[23] mux2
x4[22] i_instruction[15] net11[22] net7[22] net6 net9[22] mux2
x4[21] i_instruction[15] net11[21] net7[21] net6 net9[21] mux2
x4[20] i_instruction[15] net11[20] net7[20] net6 net9[20] mux2
x4[19] i_instruction[15] net11[19] net7[19] net6 net9[19] mux2
x4[18] i_instruction[15] net11[18] net7[18] net6 net9[18] mux2
x4[17] i_instruction[15] net11[17] net7[17] net6 net9[17] mux2
x4[16] i_instruction[15] net11[16] net7[16] net6 net9[16] mux2
x4[15] i_instruction[15] net11[15] net7[15] net6 net9[15] mux2
x4[14] i_instruction[15] net11[14] net7[14] net6 net9[14] mux2
x4[13] i_instruction[15] net11[13] net7[13] net6 net9[13] mux2
x4[12] i_instruction[15] net11[12] net7[12] net6 net9[12] mux2
x4[11] i_instruction[15] net11[11] net7[11] net6 net9[11] mux2
x4[10] i_instruction[15] net11[10] net7[10] net6 net9[10] mux2
x4[9] i_instruction[15] net11[9] net7[9] net6 net9[9] mux2
x4[8] i_instruction[15] net11[8] net7[8] net6 net9[8] mux2
x4[7] i_instruction[15] net11[7] net7[7] net6 net9[7] mux2
x4[6] i_instruction[15] net11[6] net7[6] net6 net9[6] mux2
x4[5] i_instruction[15] net11[5] net7[5] net6 net9[5] mux2
x4[4] i_instruction[15] net11[4] net7[4] net6 net9[4] mux2
x4[3] i_instruction[15] net11[3] net7[3] net6 net9[3] mux2
x4[2] i_instruction[15] net11[2] net7[2] net6 net9[2] mux2
x4[1] i_instruction[15] net11[1] net7[1] net6 net9[1] mux2
x4[0] i_instruction[15] net11[0] net7[0] net6 net9[0] mux2
x5 i_instruction[15] VSS VSS VCC VCC net6 sky130_fd_sc_hd__inv_1
x5[32] i_instruction[14] VSS net9[32] net8 net14[32] mux2
x5[31] i_instruction[14] VSS net9[31] net8 net14[31] mux2
x5[30] i_instruction[14] VSS net9[30] net8 net14[30] mux2
x5[29] i_instruction[14] VSS net9[29] net8 net14[29] mux2
x5[28] i_instruction[14] VSS net9[28] net8 net14[28] mux2
x5[27] i_instruction[14] VSS net9[27] net8 net14[27] mux2
x5[26] i_instruction[14] i_instruction[5] net9[26] net8 net14[26] mux2
x5[25] i_instruction[14] i_instruction[12] net9[25] net8 net14[25] mux2
x5[24] i_instruction[14] i_instruction[11] net9[24] net8 net14[24] mux2
x5[23] i_instruction[14] i_instruction[10] net9[23] net8 net14[23] mux2
x5[22] i_instruction[14] i_instruction[6] net9[22] net8 net14[22] mux2
x5[21] i_instruction[14] VSS net9[21] net8 net14[21] mux2
x5[20] i_instruction[14] VSS net9[20] net8 net14[20] mux2
x5[19] i_instruction[14] VSS net9[19] net8 net14[19] mux2
x5[18] i_instruction[14] VCC net9[18] net8 net14[18] mux2
x5[17] i_instruction[14] i_instruction[9] net9[17] net8 net14[17] mux2
x5[16] i_instruction[14] i_instruction[8] net9[16] net8 net14[16] mux2
x5[15] i_instruction[14] i_instruction[7] net9[15] net8 net14[15] mux2
x5[14] i_instruction[14] VSS net9[14] net8 net14[14] mux2
x5[13] i_instruction[14] VCC net9[13] net8 net14[13] mux2
x5[12] i_instruction[14] VSS net9[12] net8 net14[12] mux2
x5[11] i_instruction[14] VSS net9[11] net8 net14[11] mux2
x5[10] i_instruction[14] VCC net9[10] net8 net14[10] mux2
x5[9] i_instruction[14] i_instruction[4] net9[9] net8 net14[9] mux2
x5[8] i_instruction[14] i_instruction[3] net9[8] net8 net14[8] mux2
x5[7] i_instruction[14] i_instruction[2] net9[7] net8 net14[7] mux2
x5[6] i_instruction[14] VSS net9[6] net8 net14[6] mux2
x5[5] i_instruction[14] VSS net9[5] net8 net14[5] mux2
x5[4] i_instruction[14] VSS net9[4] net8 net14[4] mux2
x5[3] i_instruction[14] VSS net9[3] net8 net14[3] mux2
x5[2] i_instruction[14] VSS net9[2] net8 net14[2] mux2
x5[1] i_instruction[14] VCC net9[1] net8 net14[1] mux2
x5[0] i_instruction[14] VCC net9[0] net8 net14[0] mux2
x6 i_instruction[14] VSS VSS VCC VCC net8 sky130_fd_sc_hd__inv_1
x6[32] i_instruction[14] VSS net11[32] net10 VCC mux2
x6[31] i_instruction[14] VSS net11[31] net10 i_instruction[31] mux2
x6[30] i_instruction[14] VSS net11[30] net10 i_instruction[30] mux2
x6[29] i_instruction[14] VSS net11[29] net10 i_instruction[29] mux2
x6[28] i_instruction[14] VSS net11[28] net10 i_instruction[28] mux2
x6[27] i_instruction[14] VSS net11[27] net10 i_instruction[27] mux2
x6[26] i_instruction[14] i_instruction[5] net11[26] net10 i_instruction[26] mux2
x6[25] i_instruction[14] i_instruction[12] net11[25] net10 i_instruction[25] mux2
x6[24] i_instruction[14] VSS net11[24] net10 i_instruction[24] mux2
x6[23] i_instruction[14] VCC net11[23] net10 i_instruction[23] mux2
x6[22] i_instruction[14] i_instruction[4] net11[22] net10 i_instruction[22] mux2
x6[21] i_instruction[14] i_instruction[3] net11[21] net10 i_instruction[21] mux2
x6[20] i_instruction[14] i_instruction[2] net11[20] net10 i_instruction[20] mux2
x6[19] i_instruction[14] VSS net11[19] net10 i_instruction[19] mux2
x6[18] i_instruction[14] VCC net11[18] net10 i_instruction[18] mux2
x6[17] i_instruction[14] i_instruction[9] net11[17] net10 i_instruction[17] mux2
x6[16] i_instruction[14] i_instruction[8] net11[16] net10 i_instruction[16] mux2
x6[15] i_instruction[14] i_instruction[7] net11[15] net10 i_instruction[15] mux2
x6[14] i_instruction[14] VSS net11[14] net10 i_instruction[14] mux2
x6[13] i_instruction[14] VCC net11[13] net10 i_instruction[13] mux2
x6[12] i_instruction[14] VSS net11[12] net10 i_instruction[12] mux2
x6[11] i_instruction[14] i_instruction[11] net11[11] net10 i_instruction[11] mux2
x6[10] i_instruction[14] i_instruction[10] net11[10] net10 i_instruction[10] mux2
x6[9] i_instruction[14] i_instruction[6] net11[9] net10 i_instruction[9] mux2
x6[8] i_instruction[14] VSS net11[8] net10 i_instruction[8] mux2
x6[7] i_instruction[14] VSS net11[7] net10 i_instruction[7] mux2
x6[6] i_instruction[14] VSS net11[6] net10 i_instruction[6] mux2
x6[5] i_instruction[14] VCC net11[5] net10 i_instruction[5] mux2
x6[4] i_instruction[14] VSS net11[4] net10 i_instruction[4] mux2
x6[3] i_instruction[14] VSS net11[3] net10 i_instruction[3] mux2
x6[2] i_instruction[14] VSS net11[2] net10 i_instruction[2] mux2
x6[1] i_instruction[14] VCC net11[1] net10 i_instruction[1] mux2
x6[0] i_instruction[14] VCC net11[0] net10 i_instruction[0] mux2
x7 i_instruction[14] VSS VSS VCC VCC net10 sky130_fd_sc_hd__inv_1
x7[32] net12 VSS net14[32] net13 VSS mux2
x7[31] net12 VSS net14[31] net13 VSS mux2
x7[30] net12 VSS net14[30] net13 VSS mux2
x7[29] net12 i_instruction[10] net14[29] net13 VSS mux2
x7[28] net12 i_instruction[9] net14[28] net13 VSS mux2
x7[27] net12 i_instruction[8] net14[27] net13 VSS mux2
x7[26] net12 i_instruction[7] net14[26] net13 VSS mux2
x7[25] net12 i_instruction[12] net14[25] net13 VSS mux2
x7[24] net12 i_instruction[11] net14[24] net13 VSS mux2
x7[23] net12 i_instruction[5] net14[23] net13 VSS mux2
x7[22] net12 i_instruction[6] net14[22] net13 VSS mux2
x7[21] net12 VSS net14[21] net13 VSS mux2
x7[20] net12 VSS net14[20] net13 VSS mux2
x7[19] net12 VSS net14[19] net13 VSS mux2
x7[18] net12 VSS net14[18] net13 VSS mux2
x7[17] net12 VSS net14[17] net13 VSS mux2
x7[16] net12 VCC net14[16] net13 VSS mux2
x7[15] net12 VSS net14[15] net13 VSS mux2
x7[14] net12 VSS net14[14] net13 VSS mux2
x7[13] net12 VSS net14[13] net13 VSS mux2
x7[12] net12 VSS net14[12] net13 VSS mux2
x7[11] net12 VSS net14[11] net13 VSS mux2
x7[10] net12 VCC net14[10] net13 VSS mux2
x7[9] net12 i_instruction[4] net14[9] net13 VSS mux2
x7[8] net12 i_instruction[3] net14[8] net13 VSS mux2
x7[7] net12 i_instruction[2] net14[7] net13 VSS mux2
x7[6] net12 VSS net14[6] net13 VSS mux2
x7[5] net12 VSS net14[5] net13 VSS mux2
x7[4] net12 VCC net14[4] net13 VSS mux2
x7[3] net12 VSS net14[3] net13 VSS mux2
x7[2] net12 VSS net14[2] net13 VSS mux2
x7[1] net12 VCC net14[1] net13 VSS mux2
x7[0] net12 VCC net14[0] net13 VSS mux2
x8 net12 VSS VSS VCC VCC net13 sky130_fd_sc_hd__inv_1
x2 i_instruction[12] i_instruction[11] i_instruction[10] VSS VSS VCC VCC net15
+ sky130_fd_sc_hd__or3_1
x9 i_instruction[9] i_instruction[8] i_instruction[7] VSS VSS VCC VCC net61 sky130_fd_sc_hd__or3_1
x10 i_instruction[6] i_instruction[5] VSS VSS VCC VCC net16 sky130_fd_sc_hd__or2_1
x11 net15 net61 net16 VSS VSS VCC VCC net12 sky130_fd_sc_hd__or3_1
x8[32] i_instruction[15] net22[32] net18[32] net17 net21[32] mux2
x8[31] i_instruction[15] net22[31] net18[31] net17 net21[31] mux2
x8[30] i_instruction[15] net22[30] net18[30] net17 net21[30] mux2
x8[29] i_instruction[15] net22[29] net18[29] net17 net21[29] mux2
x8[28] i_instruction[15] net22[28] net18[28] net17 net21[28] mux2
x8[27] i_instruction[15] net22[27] net18[27] net17 net21[27] mux2
x8[26] i_instruction[15] net22[26] net18[26] net17 net21[26] mux2
x8[25] i_instruction[15] net22[25] net18[25] net17 net21[25] mux2
x8[24] i_instruction[15] net22[24] net18[24] net17 net21[24] mux2
x8[23] i_instruction[15] net22[23] net18[23] net17 net21[23] mux2
x8[22] i_instruction[15] net22[22] net18[22] net17 net21[22] mux2
x8[21] i_instruction[15] net22[21] net18[21] net17 net21[21] mux2
x8[20] i_instruction[15] net22[20] net18[20] net17 net21[20] mux2
x8[19] i_instruction[15] net22[19] net18[19] net17 net21[19] mux2
x8[18] i_instruction[15] net22[18] net18[18] net17 net21[18] mux2
x8[17] i_instruction[15] net22[17] net18[17] net17 net21[17] mux2
x8[16] i_instruction[15] net22[16] net18[16] net17 net21[16] mux2
x8[15] i_instruction[15] net22[15] net18[15] net17 net21[15] mux2
x8[14] i_instruction[15] net22[14] net18[14] net17 net21[14] mux2
x8[13] i_instruction[15] net22[13] net18[13] net17 net21[13] mux2
x8[12] i_instruction[15] net22[12] net18[12] net17 net21[12] mux2
x8[11] i_instruction[15] net22[11] net18[11] net17 net21[11] mux2
x8[10] i_instruction[15] net22[10] net18[10] net17 net21[10] mux2
x8[9] i_instruction[15] net22[9] net18[9] net17 net21[9] mux2
x8[8] i_instruction[15] net22[8] net18[8] net17 net21[8] mux2
x8[7] i_instruction[15] net22[7] net18[7] net17 net21[7] mux2
x8[6] i_instruction[15] net22[6] net18[6] net17 net21[6] mux2
x8[5] i_instruction[15] net22[5] net18[5] net17 net21[5] mux2
x8[4] i_instruction[15] net22[4] net18[4] net17 net21[4] mux2
x8[3] i_instruction[15] net22[3] net18[3] net17 net21[3] mux2
x8[2] i_instruction[15] net22[2] net18[2] net17 net21[2] mux2
x8[1] i_instruction[15] net22[1] net18[1] net17 net21[1] mux2
x8[0] i_instruction[15] net22[0] net18[0] net17 net21[0] mux2
x12 i_instruction[15] VSS VSS VCC VCC net17 sky130_fd_sc_hd__inv_1
x9[32] i_instruction[14] VSS net22[32] net19 net48[32] mux2
x9[31] i_instruction[14] i_instruction[12] net22[31] net19 net48[31] mux2
x9[30] i_instruction[14] i_instruction[12] net22[30] net19 net48[30] mux2
x9[29] i_instruction[14] i_instruction[12] net22[29] net19 net48[29] mux2
x9[28] i_instruction[14] i_instruction[12] net22[28] net19 net48[28] mux2
x9[27] i_instruction[14] i_instruction[6] net22[27] net19 net48[27] mux2
x9[26] i_instruction[14] i_instruction[5] net22[26] net19 net48[26] mux2
x9[25] i_instruction[14] i_instruction[2] net22[25] net19 net48[25] mux2
x9[24] i_instruction[14] VSS net22[24] net19 net48[24] mux2
x9[23] i_instruction[14] VSS net22[23] net19 net48[23] mux2
x9[22] i_instruction[14] VSS net22[22] net19 net48[22] mux2
x9[21] i_instruction[14] VSS net22[21] net19 net48[21] mux2
x9[20] i_instruction[14] VSS net22[20] net19 net48[20] mux2
x9[19] i_instruction[14] VSS net22[19] net19 net48[19] mux2
x9[18] i_instruction[14] VCC net22[18] net19 net48[18] mux2
x9[17] i_instruction[14] i_instruction[9] net22[17] net19 net48[17] mux2
x9[16] i_instruction[14] i_instruction[8] net22[16] net19 net48[16] mux2
x9[15] i_instruction[14] i_instruction[7] net22[15] net19 net48[15] mux2
x9[14] i_instruction[14] VSS net22[14] net19 net48[14] mux2
x9[13] i_instruction[14] VSS net22[13] net19 net48[13] mux2
x9[12] i_instruction[14] i_instruction[13] net22[12] net19 net48[12] mux2
x9[11] i_instruction[14] i_instruction[11] net22[11] net19 net48[11] mux2
x9[10] i_instruction[14] i_instruction[10] net22[10] net19 net48[10] mux2
x9[9] i_instruction[14] i_instruction[4] net22[9] net19 net48[9] mux2
x9[8] i_instruction[14] i_instruction[3] net22[8] net19 net48[8] mux2
x9[7] i_instruction[14] i_instruction[12] net22[7] net19 net48[7] mux2
x9[6] i_instruction[14] VCC net22[6] net19 net48[6] mux2
x9[5] i_instruction[14] VCC net22[5] net19 net48[5] mux2
x9[4] i_instruction[14] VSS net22[4] net19 net48[4] mux2
x9[3] i_instruction[14] VSS net22[3] net19 net48[3] mux2
x9[2] i_instruction[14] VSS net22[2] net19 net48[2] mux2
x9[1] i_instruction[14] VCC net22[1] net19 net48[1] mux2
x9[0] i_instruction[14] VCC net22[0] net19 net48[0] mux2
x13 i_instruction[14] VSS VSS VCC VCC net19 sky130_fd_sc_hd__inv_1
x10[32] i_instruction[14] net27[32] net21[32] net20 net26[32] mux2
x10[31] i_instruction[14] net27[31] net21[31] net20 net26[31] mux2
x10[30] i_instruction[14] net27[30] net21[30] net20 net26[30] mux2
x10[29] i_instruction[14] net27[29] net21[29] net20 net26[29] mux2
x10[28] i_instruction[14] net27[28] net21[28] net20 net26[28] mux2
x10[27] i_instruction[14] net27[27] net21[27] net20 net26[27] mux2
x10[26] i_instruction[14] net27[26] net21[26] net20 net26[26] mux2
x10[25] i_instruction[14] net27[25] net21[25] net20 net26[25] mux2
x10[24] i_instruction[14] net27[24] net21[24] net20 net26[24] mux2
x10[23] i_instruction[14] net27[23] net21[23] net20 net26[23] mux2
x10[22] i_instruction[14] net27[22] net21[22] net20 net26[22] mux2
x10[21] i_instruction[14] net27[21] net21[21] net20 net26[21] mux2
x10[20] i_instruction[14] net27[20] net21[20] net20 net26[20] mux2
x10[19] i_instruction[14] net27[19] net21[19] net20 net26[19] mux2
x10[18] i_instruction[14] net27[18] net21[18] net20 net26[18] mux2
x10[17] i_instruction[14] net27[17] net21[17] net20 net26[17] mux2
x10[16] i_instruction[14] net27[16] net21[16] net20 net26[16] mux2
x10[15] i_instruction[14] net27[15] net21[15] net20 net26[15] mux2
x10[14] i_instruction[14] net27[14] net21[14] net20 net26[14] mux2
x10[13] i_instruction[14] net27[13] net21[13] net20 net26[13] mux2
x10[12] i_instruction[14] net27[12] net21[12] net20 net26[12] mux2
x10[11] i_instruction[14] net27[11] net21[11] net20 net26[11] mux2
x10[10] i_instruction[14] net27[10] net21[10] net20 net26[10] mux2
x10[9] i_instruction[14] net27[9] net21[9] net20 net26[9] mux2
x10[8] i_instruction[14] net27[8] net21[8] net20 net26[8] mux2
x10[7] i_instruction[14] net27[7] net21[7] net20 net26[7] mux2
x10[6] i_instruction[14] net27[6] net21[6] net20 net26[6] mux2
x10[5] i_instruction[14] net27[5] net21[5] net20 net26[5] mux2
x10[4] i_instruction[14] net27[4] net21[4] net20 net26[4] mux2
x10[3] i_instruction[14] net27[3] net21[3] net20 net26[3] mux2
x10[2] i_instruction[14] net27[2] net21[2] net20 net26[2] mux2
x10[1] i_instruction[14] net27[1] net21[1] net20 net26[1] mux2
x10[0] i_instruction[14] net27[0] net21[0] net20 net26[0] mux2
x14 i_instruction[14] VSS VSS VCC VCC net20 sky130_fd_sc_hd__inv_1
x11[32] i_instruction[13] VSS net26[32] net23 VSS mux2
x11[31] i_instruction[13] i_instruction[12] net26[31] net23 i_instruction[12] mux2
x11[30] i_instruction[13] i_instruction[8] net26[30] net23 i_instruction[12] mux2
x11[29] i_instruction[13] i_instruction[10] net26[29] net23 i_instruction[12] mux2
x11[28] i_instruction[13] i_instruction[9] net26[28] net23 i_instruction[12] mux2
x11[27] i_instruction[13] i_instruction[6] net26[27] net23 i_instruction[12] mux2
x11[26] i_instruction[13] i_instruction[7] net26[26] net23 i_instruction[12] mux2
x11[25] i_instruction[13] i_instruction[2] net26[25] net23 i_instruction[12] mux2
x11[24] i_instruction[13] i_instruction[11] net26[24] net23 i_instruction[6] mux2
x11[23] i_instruction[13] i_instruction[5] net26[23] net23 i_instruction[5] mux2
x11[22] i_instruction[13] i_instruction[4] net26[22] net23 i_instruction[4] mux2
x11[21] i_instruction[13] i_instruction[3] net26[21] net23 i_instruction[3] mux2
x11[20] i_instruction[13] i_instruction[12] net26[20] net23 i_instruction[2] mux2
x11[19] i_instruction[13] i_instruction[12] net26[19] net23 i_instruction[11] mux2
x11[18] i_instruction[13] i_instruction[12] net26[18] net23 i_instruction[10] mux2
x11[17] i_instruction[13] i_instruction[12] net26[17] net23 i_instruction[9] mux2
x11[16] i_instruction[13] i_instruction[12] net26[16] net23 i_instruction[8] mux2
x11[15] i_instruction[13] i_instruction[12] net26[15] net23 i_instruction[7] mux2
x11[14] i_instruction[13] i_instruction[12] net26[14] net23 VSS mux2
x11[13] i_instruction[13] i_instruction[12] net26[13] net23 VSS mux2
x11[12] i_instruction[13] i_instruction[12] net26[12] net23 VSS mux2
x11[11] i_instruction[13] VSS net26[11] net23 i_instruction[11] mux2
x11[10] i_instruction[13] VSS net26[10] net23 i_instruction[10] mux2
x11[9] i_instruction[13] VSS net26[9] net23 i_instruction[9] mux2
x11[8] i_instruction[13] VSS net26[8] net23 i_instruction[8] mux2
x11[7] i_instruction[13] VCC net26[7] net23 i_instruction[7] mux2
x11[6] i_instruction[13] VCC net26[6] net23 VSS mux2
x11[5] i_instruction[13] VCC net26[5] net23 VSS mux2
x11[4] i_instruction[13] VSS net26[4] net23 VCC mux2
x11[3] i_instruction[13] VCC net26[3] net23 VSS mux2
x11[2] i_instruction[13] VCC net26[2] net23 VSS mux2
x11[1] i_instruction[13] VCC net26[1] net23 VCC mux2
x11[0] i_instruction[13] VCC net26[0] net23 VCC mux2
x15 i_instruction[13] VSS VSS VCC VCC net23 sky130_fd_sc_hd__inv_1
x12[32] i_instruction[13] net30[32] net27[32] net24 VSS mux2
x12[31] i_instruction[13] net30[31] net27[31] net24 i_instruction[12] mux2
x12[30] i_instruction[13] net30[30] net27[30] net24 i_instruction[12] mux2
x12[29] i_instruction[13] net30[29] net27[29] net24 i_instruction[12] mux2
x12[28] i_instruction[13] net30[28] net27[28] net24 i_instruction[12] mux2
x12[27] i_instruction[13] net30[27] net27[27] net24 i_instruction[12] mux2
x12[26] i_instruction[13] net30[26] net27[26] net24 i_instruction[12] mux2
x12[25] i_instruction[13] net30[25] net27[25] net24 i_instruction[12] mux2
x12[24] i_instruction[13] net30[24] net27[24] net24 i_instruction[6] mux2
x12[23] i_instruction[13] net30[23] net27[23] net24 i_instruction[5] mux2
x12[22] i_instruction[13] net30[22] net27[22] net24 i_instruction[4] mux2
x12[21] i_instruction[13] net30[21] net27[21] net24 i_instruction[3] mux2
x12[20] i_instruction[13] net30[20] net27[20] net24 i_instruction[2] mux2
x12[19] i_instruction[13] net30[19] net27[19] net24 VSS mux2
x12[18] i_instruction[13] net30[18] net27[18] net24 VSS mux2
x12[17] i_instruction[13] net30[17] net27[17] net24 VSS mux2
x12[16] i_instruction[13] net30[16] net27[16] net24 VSS mux2
x12[15] i_instruction[13] net30[15] net27[15] net24 VSS mux2
x12[14] i_instruction[13] net30[14] net27[14] net24 VSS mux2
x12[13] i_instruction[13] net30[13] net27[13] net24 VSS mux2
x12[12] i_instruction[13] net30[12] net27[12] net24 VSS mux2
x12[11] i_instruction[13] net30[11] net27[11] net24 i_instruction[11] mux2
x12[10] i_instruction[13] net30[10] net27[10] net24 i_instruction[10] mux2
x12[9] i_instruction[13] net30[9] net27[9] net24 i_instruction[9] mux2
x12[8] i_instruction[13] net30[8] net27[8] net24 i_instruction[8] mux2
x12[7] i_instruction[13] net30[7] net27[7] net24 i_instruction[7] mux2
x12[6] i_instruction[13] net30[6] net27[6] net24 VSS mux2
x12[5] i_instruction[13] net30[5] net27[5] net24 VSS mux2
x12[4] i_instruction[13] net30[4] net27[4] net24 VCC mux2
x12[3] i_instruction[13] net30[3] net27[3] net24 VSS mux2
x12[2] i_instruction[13] net30[2] net27[2] net24 VSS mux2
x12[1] i_instruction[13] net30[1] net27[1] net24 VCC mux2
x12[0] i_instruction[13] net30[0] net27[0] net24 VCC mux2
x16 i_instruction[13] VSS VSS VCC VCC net24 sky130_fd_sc_hd__inv_1
x13[32] i_instruction[13] VSS net48[32] net25 net34[32] mux2
x13[31] i_instruction[13] i_instruction[12] net48[31] net25 net34[31] mux2
x13[30] i_instruction[13] i_instruction[8] net48[30] net25 net34[30] mux2
x13[29] i_instruction[13] i_instruction[10] net48[29] net25 net34[29] mux2
x13[28] i_instruction[13] i_instruction[9] net48[28] net25 net34[28] mux2
x13[27] i_instruction[13] i_instruction[6] net48[27] net25 net34[27] mux2
x13[26] i_instruction[13] i_instruction[7] net48[26] net25 net34[26] mux2
x13[25] i_instruction[13] i_instruction[2] net48[25] net25 net34[25] mux2
x13[24] i_instruction[13] i_instruction[11] net48[24] net25 net34[24] mux2
x13[23] i_instruction[13] i_instruction[5] net48[23] net25 net34[23] mux2
x13[22] i_instruction[13] i_instruction[4] net48[22] net25 net34[22] mux2
x13[21] i_instruction[13] i_instruction[3] net48[21] net25 net34[21] mux2
x13[20] i_instruction[13] i_instruction[12] net48[20] net25 net34[20] mux2
x13[19] i_instruction[13] i_instruction[12] net48[19] net25 net34[19] mux2
x13[18] i_instruction[13] i_instruction[12] net48[18] net25 net34[18] mux2
x13[17] i_instruction[13] i_instruction[12] net48[17] net25 net34[17] mux2
x13[16] i_instruction[13] i_instruction[12] net48[16] net25 net34[16] mux2
x13[15] i_instruction[13] i_instruction[12] net48[15] net25 net34[15] mux2
x13[14] i_instruction[13] i_instruction[12] net48[14] net25 net34[14] mux2
x13[13] i_instruction[13] i_instruction[12] net48[13] net25 net34[13] mux2
x13[12] i_instruction[13] i_instruction[12] net48[12] net25 net34[12] mux2
x13[11] i_instruction[13] VSS net48[11] net25 net34[11] mux2
x13[10] i_instruction[13] VSS net48[10] net25 net34[10] mux2
x13[9] i_instruction[13] VSS net48[9] net25 net34[9] mux2
x13[8] i_instruction[13] VSS net48[8] net25 net34[8] mux2
x13[7] i_instruction[13] VSS net48[7] net25 net34[7] mux2
x13[6] i_instruction[13] VCC net48[6] net25 net34[6] mux2
x13[5] i_instruction[13] VCC net48[5] net25 net34[5] mux2
x13[4] i_instruction[13] VSS net48[4] net25 net34[4] mux2
x13[3] i_instruction[13] VCC net48[3] net25 net34[3] mux2
x13[2] i_instruction[13] VCC net48[2] net25 net34[2] mux2
x13[1] i_instruction[13] VCC net48[1] net25 net34[1] mux2
x13[0] i_instruction[13] VCC net48[0] net25 net34[0] mux2
x17 i_instruction[13] VSS VSS VCC VCC net25 sky130_fd_sc_hd__inv_1
x15[32] net29 VSS net30[32] net28 VSS mux2
x15[31] net29 i_instruction[12] net30[31] net28 i_instruction[12] mux2
x15[30] net29 i_instruction[12] net30[30] net28 i_instruction[12] mux2
x15[29] net29 i_instruction[12] net30[29] net28 i_instruction[12] mux2
x15[28] net29 i_instruction[4] net30[28] net28 i_instruction[12] mux2
x15[27] net29 i_instruction[3] net30[27] net28 i_instruction[12] mux2
x15[26] net29 i_instruction[5] net30[26] net28 i_instruction[12] mux2
x15[25] net29 i_instruction[2] net30[25] net28 i_instruction[12] mux2
x15[24] net29 i_instruction[6] net30[24] net28 i_instruction[12] mux2
x15[23] net29 VSS net30[23] net28 i_instruction[12] mux2
x15[22] net29 VSS net30[22] net28 i_instruction[12] mux2
x15[21] net29 VSS net30[21] net28 i_instruction[12] mux2
x15[20] net29 VSS net30[20] net28 i_instruction[12] mux2
x15[19] net29 VSS net30[19] net28 i_instruction[12] mux2
x15[18] net29 VSS net30[18] net28 i_instruction[12] mux2
x15[17] net29 VSS net30[17] net28 i_instruction[12] mux2
x15[16] net29 VCC net30[16] net28 i_instruction[6] mux2
x15[15] net29 VSS net30[15] net28 i_instruction[5] mux2
x15[14] net29 VSS net30[14] net28 i_instruction[4] mux2
x15[13] net29 VSS net30[13] net28 i_instruction[3] mux2
x15[12] net29 VSS net30[12] net28 i_instruction[2] mux2
x15[11] net29 VSS net30[11] net28 i_instruction[11] mux2
x15[10] net29 VSS net30[10] net28 i_instruction[10] mux2
x15[9] net29 VSS net30[9] net28 i_instruction[9] mux2
x15[8] net29 VCC net30[8] net28 i_instruction[8] mux2
x15[7] net29 VSS net30[7] net28 i_instruction[7] mux2
x15[6] net29 VSS net30[6] net28 VSS mux2
x15[5] net29 VSS net30[5] net28 VCC mux2
x15[4] net29 VCC net30[4] net28 VCC mux2
x15[3] net29 VSS net30[3] net28 VSS mux2
x15[2] net29 VSS net30[2] net28 VCC mux2
x15[1] net29 VCC net30[1] net28 VCC mux2
x15[0] net29 VCC net30[0] net28 VCC mux2
x20 net29 VSS VSS VCC VCC net28 sky130_fd_sc_hd__inv_1
x21 net62 net63 net64 VSS VSS VCC VCC net65 sky130_fd_sc_hd__and3_1
x22 i_instruction[8] net66 VSS VSS VCC VCC net31 sky130_fd_sc_hd__and2_1
x23 net65 net31 VSS VSS VCC VCC net29 sky130_fd_sc_hd__and2_1
x24 i_instruction[11] VSS VSS VCC VCC net62 sky130_fd_sc_hd__inv_1
x25 i_instruction[10] VSS VSS VCC VCC net63 sky130_fd_sc_hd__inv_1
x26 i_instruction[9] VSS VSS VCC VCC net64 sky130_fd_sc_hd__inv_1
x27 i_instruction[7] VSS VSS VCC VCC net66 sky130_fd_sc_hd__inv_1
x14[32] i_instruction[11] net35[32] net34[32] net32 VSS mux2
x14[31] i_instruction[11] net35[31] net34[31] net32 VSS mux2
x14[30] i_instruction[11] net35[30] net34[30] net32 i_instruction[10] mux2
x14[29] i_instruction[11] net35[29] net34[29] net32 VSS mux2
x14[28] i_instruction[11] net35[28] net34[28] net32 VSS mux2
x14[27] i_instruction[11] net35[27] net34[27] net32 VSS mux2
x14[26] i_instruction[11] net35[26] net34[26] net32 VSS mux2
x14[25] i_instruction[11] net35[25] net34[25] net32 VSS mux2
x14[24] i_instruction[11] net35[24] net34[24] net32 i_instruction[6] mux2
x14[23] i_instruction[11] net35[23] net34[23] net32 i_instruction[5] mux2
x14[22] i_instruction[11] net35[22] net34[22] net32 i_instruction[4] mux2
x14[21] i_instruction[11] net35[21] net34[21] net32 i_instruction[3] mux2
x14[20] i_instruction[11] net35[20] net34[20] net32 i_instruction[2] mux2
x14[19] i_instruction[11] net35[19] net34[19] net32 VSS mux2
x14[18] i_instruction[11] net35[18] net34[18] net32 VCC mux2
x14[17] i_instruction[11] net35[17] net34[17] net32 i_instruction[9] mux2
x14[16] i_instruction[11] net35[16] net34[16] net32 i_instruction[8] mux2
x14[15] i_instruction[11] net35[15] net34[15] net32 i_instruction[7] mux2
x14[14] i_instruction[11] net35[14] net34[14] net32 VCC mux2
x14[13] i_instruction[11] net35[13] net34[13] net32 VSS mux2
x14[12] i_instruction[11] net35[12] net34[12] net32 VCC mux2
x14[11] i_instruction[11] net35[11] net34[11] net32 VSS mux2
x14[10] i_instruction[11] net35[10] net34[10] net32 VCC mux2
x14[9] i_instruction[11] net35[9] net34[9] net32 i_instruction[9] mux2
x14[8] i_instruction[11] net35[8] net34[8] net32 i_instruction[8] mux2
x14[7] i_instruction[11] net35[7] net34[7] net32 i_instruction[7] mux2
x14[6] i_instruction[11] net35[6] net34[6] net32 VSS mux2
x14[5] i_instruction[11] net35[5] net34[5] net32 VSS mux2
x14[4] i_instruction[11] net35[4] net34[4] net32 VCC mux2
x14[3] i_instruction[11] net35[3] net34[3] net32 VSS mux2
x14[2] i_instruction[11] net35[2] net34[2] net32 VSS mux2
x14[1] i_instruction[11] net35[1] net34[1] net32 VCC mux2
x14[0] i_instruction[11] net35[0] net34[0] net32 VCC mux2
x18 i_instruction[11] VSS VSS VCC VCC net32 sky130_fd_sc_hd__inv_1
x17[32] i_instruction[10] net41[32] net35[32] net33 VSS mux2
x17[31] i_instruction[10] net41[31] net35[31] net33 i_instruction[12] mux2
x17[30] i_instruction[10] net41[30] net35[30] net33 i_instruction[12] mux2
x17[29] i_instruction[10] net41[29] net35[29] net33 i_instruction[12] mux2
x17[28] i_instruction[10] net41[28] net35[28] net33 i_instruction[12] mux2
x17[27] i_instruction[10] net41[27] net35[27] net33 i_instruction[12] mux2
x17[26] i_instruction[10] net41[26] net35[26] net33 i_instruction[12] mux2
x17[25] i_instruction[10] net41[25] net35[25] net33 i_instruction[12] mux2
x17[24] i_instruction[10] net41[24] net35[24] net33 i_instruction[6] mux2
x17[23] i_instruction[10] net41[23] net35[23] net33 i_instruction[5] mux2
x17[22] i_instruction[10] net41[22] net35[22] net33 i_instruction[4] mux2
x17[21] i_instruction[10] net41[21] net35[21] net33 i_instruction[3] mux2
x17[20] i_instruction[10] net41[20] net35[20] net33 i_instruction[2] mux2
x17[19] i_instruction[10] net41[19] net35[19] net33 VSS mux2
x17[18] i_instruction[10] net41[18] net35[18] net33 VCC mux2
x17[17] i_instruction[10] net41[17] net35[17] net33 i_instruction[9] mux2
x17[16] i_instruction[10] net41[16] net35[16] net33 i_instruction[8] mux2
x17[15] i_instruction[10] net41[15] net35[15] net33 i_instruction[7] mux2
x17[14] i_instruction[10] net41[14] net35[14] net33 VCC mux2
x17[13] i_instruction[10] net41[13] net35[13] net33 VCC mux2
x17[12] i_instruction[10] net41[12] net35[12] net33 VCC mux2
x17[11] i_instruction[10] net41[11] net35[11] net33 VSS mux2
x17[10] i_instruction[10] net41[10] net35[10] net33 VCC mux2
x17[9] i_instruction[10] net41[9] net35[9] net33 i_instruction[9] mux2
x17[8] i_instruction[10] net41[8] net35[8] net33 i_instruction[8] mux2
x17[7] i_instruction[10] net41[7] net35[7] net33 i_instruction[7] mux2
x17[6] i_instruction[10] net41[6] net35[6] net33 VSS mux2
x17[5] i_instruction[10] net41[5] net35[5] net33 VSS mux2
x17[4] i_instruction[10] net41[4] net35[4] net33 VCC mux2
x17[3] i_instruction[10] net41[3] net35[3] net33 VSS mux2
x17[2] i_instruction[10] net41[2] net35[2] net33 VSS mux2
x17[1] i_instruction[10] net41[1] net35[1] net33 VCC mux2
x17[0] i_instruction[10] net41[0] net35[0] net33 VCC mux2
x28 i_instruction[10] VSS VSS VCC VCC net33 sky130_fd_sc_hd__inv_1
x16[32] i_instruction[6] net40[32] net41[32] net36 net39[32] mux2
x16[31] i_instruction[6] net40[31] net41[31] net36 net39[31] mux2
x16[30] i_instruction[6] net40[30] net41[30] net36 net39[30] mux2
x16[29] i_instruction[6] net40[29] net41[29] net36 net39[29] mux2
x16[28] i_instruction[6] net40[28] net41[28] net36 net39[28] mux2
x16[27] i_instruction[6] net40[27] net41[27] net36 net39[27] mux2
x16[26] i_instruction[6] net40[26] net41[26] net36 net39[26] mux2
x16[25] i_instruction[6] net40[25] net41[25] net36 net39[25] mux2
x16[24] i_instruction[6] net40[24] net41[24] net36 net39[24] mux2
x16[23] i_instruction[6] net40[23] net41[23] net36 net39[23] mux2
x16[22] i_instruction[6] net40[22] net41[22] net36 net39[22] mux2
x16[21] i_instruction[6] net40[21] net41[21] net36 net39[21] mux2
x16[20] i_instruction[6] net40[20] net41[20] net36 net39[20] mux2
x16[19] i_instruction[6] net40[19] net41[19] net36 net39[19] mux2
x16[18] i_instruction[6] net40[18] net41[18] net36 net39[18] mux2
x16[17] i_instruction[6] net40[17] net41[17] net36 net39[17] mux2
x16[16] i_instruction[6] net40[16] net41[16] net36 net39[16] mux2
x16[15] i_instruction[6] net40[15] net41[15] net36 net39[15] mux2
x16[14] i_instruction[6] net40[14] net41[14] net36 net39[14] mux2
x16[13] i_instruction[6] net40[13] net41[13] net36 net39[13] mux2
x16[12] i_instruction[6] net40[12] net41[12] net36 net39[12] mux2
x16[11] i_instruction[6] net40[11] net41[11] net36 net39[11] mux2
x16[10] i_instruction[6] net40[10] net41[10] net36 net39[10] mux2
x16[9] i_instruction[6] net40[9] net41[9] net36 net39[9] mux2
x16[8] i_instruction[6] net40[8] net41[8] net36 net39[8] mux2
x16[7] i_instruction[6] net40[7] net41[7] net36 net39[7] mux2
x16[6] i_instruction[6] net40[6] net41[6] net36 net39[6] mux2
x16[5] i_instruction[6] net40[5] net41[5] net36 net39[5] mux2
x16[4] i_instruction[6] net40[4] net41[4] net36 net39[4] mux2
x16[3] i_instruction[6] net40[3] net41[3] net36 net39[3] mux2
x16[2] i_instruction[6] net40[2] net41[2] net36 net39[2] mux2
x16[1] i_instruction[6] net40[1] net41[1] net36 net39[1] mux2
x16[0] i_instruction[6] net40[0] net41[0] net36 net39[0] mux2
x19 i_instruction[6] VSS VSS VCC VCC net36 sky130_fd_sc_hd__inv_1
x18[32] i_instruction[5] VSS net39[32] net37 VSS mux2
x18[31] i_instruction[5] VSS net39[31] net37 VSS mux2
x18[30] i_instruction[5] VSS net39[30] net37 VCC mux2
x18[29] i_instruction[5] VSS net39[29] net37 VSS mux2
x18[28] i_instruction[5] VSS net39[28] net37 VSS mux2
x18[27] i_instruction[5] VSS net39[27] net37 VSS mux2
x18[26] i_instruction[5] VSS net39[26] net37 VSS mux2
x18[25] i_instruction[5] VSS net39[25] net37 VSS mux2
x18[24] i_instruction[5] VSS net39[24] net37 VSS mux2
x18[23] i_instruction[5] VCC net39[23] net37 VCC mux2
x18[22] i_instruction[5] i_instruction[4] net39[22] net37 i_instruction[4] mux2
x18[21] i_instruction[5] i_instruction[3] net39[21] net37 i_instruction[3] mux2
x18[20] i_instruction[5] i_instruction[2] net39[20] net37 i_instruction[2] mux2
x18[19] i_instruction[5] VSS net39[19] net37 VSS mux2
x18[18] i_instruction[5] VCC net39[18] net37 VCC mux2
x18[17] i_instruction[5] i_instruction[9] net39[17] net37 i_instruction[9] mux2
x18[16] i_instruction[5] i_instruction[8] net39[16] net37 i_instruction[8] mux2
x18[15] i_instruction[5] i_instruction[7] net39[15] net37 i_instruction[7] mux2
x18[14] i_instruction[5] VCC net39[14] net37 VSS mux2
x18[13] i_instruction[5] VSS net39[13] net37 VSS mux2
x18[12] i_instruction[5] VSS net39[12] net37 VSS mux2
x18[11] i_instruction[5] VSS net39[11] net37 VSS mux2
x18[10] i_instruction[5] VCC net39[10] net37 VCC mux2
x18[9] i_instruction[5] i_instruction[9] net39[9] net37 i_instruction[9] mux2
x18[8] i_instruction[5] i_instruction[8] net39[8] net37 i_instruction[8] mux2
x18[7] i_instruction[5] i_instruction[7] net39[7] net37 i_instruction[7] mux2
x18[6] i_instruction[5] VSS net39[6] net37 VSS mux2
x18[5] i_instruction[5] VCC net39[5] net37 VCC mux2
x18[4] i_instruction[5] VCC net39[4] net37 VCC mux2
x18[3] i_instruction[5] VSS net39[3] net37 VSS mux2
x18[2] i_instruction[5] VSS net39[2] net37 VSS mux2
x18[1] i_instruction[5] VCC net39[1] net37 VCC mux2
x18[0] i_instruction[5] VCC net39[0] net37 VCC mux2
x29 i_instruction[5] VSS VSS VCC VCC net37 sky130_fd_sc_hd__inv_1
x19[32] i_instruction[5] VSS net40[32] net38 VSS mux2
x19[31] i_instruction[5] VSS net40[31] net38 VSS mux2
x19[30] i_instruction[5] VSS net40[30] net38 VSS mux2
x19[29] i_instruction[5] VSS net40[29] net38 VSS mux2
x19[28] i_instruction[5] VSS net40[28] net38 VSS mux2
x19[27] i_instruction[5] VSS net40[27] net38 VSS mux2
x19[26] i_instruction[5] VSS net40[26] net38 VSS mux2
x19[25] i_instruction[5] VSS net40[25] net38 VSS mux2
x19[24] i_instruction[5] VSS net40[24] net38 VSS mux2
x19[23] i_instruction[5] VCC net40[23] net38 VCC mux2
x19[22] i_instruction[5] i_instruction[4] net40[22] net38 i_instruction[4] mux2
x19[21] i_instruction[5] i_instruction[3] net40[21] net38 i_instruction[3] mux2
x19[20] i_instruction[5] i_instruction[2] net40[20] net38 i_instruction[2] mux2
x19[19] i_instruction[5] VSS net40[19] net38 VSS mux2
x19[18] i_instruction[5] VCC net40[18] net38 VCC mux2
x19[17] i_instruction[5] i_instruction[9] net40[17] net38 i_instruction[9] mux2
x19[16] i_instruction[5] i_instruction[8] net40[16] net38 i_instruction[8] mux2
x19[15] i_instruction[5] i_instruction[7] net40[15] net38 i_instruction[7] mux2
x19[14] i_instruction[5] VCC net40[14] net38 VCC mux2
x19[13] i_instruction[5] VCC net40[13] net38 VCC mux2
x19[12] i_instruction[5] VCC net40[12] net38 VSS mux2
x19[11] i_instruction[5] VSS net40[11] net38 VSS mux2
x19[10] i_instruction[5] VCC net40[10] net38 VCC mux2
x19[9] i_instruction[5] i_instruction[9] net40[9] net38 i_instruction[9] mux2
x19[8] i_instruction[5] i_instruction[8] net40[8] net38 i_instruction[8] mux2
x19[7] i_instruction[5] i_instruction[7] net40[7] net38 i_instruction[7] mux2
x19[6] i_instruction[5] VSS net40[6] net38 VSS mux2
x19[5] i_instruction[5] VCC net40[5] net38 VCC mux2
x19[4] i_instruction[5] VCC net40[4] net38 VCC mux2
x19[3] i_instruction[5] VSS net40[3] net38 VSS mux2
x19[2] i_instruction[5] VSS net40[2] net38 VSS mux2
x19[1] i_instruction[5] VCC net40[1] net38 VCC mux2
x19[0] i_instruction[5] VCC net40[0] net38 VCC mux2
x30 i_instruction[5] VSS VSS VCC VCC net38 sky130_fd_sc_hd__inv_1
x20[32] i_instruction[15] net46[32] net47[32] net42 net45[32] mux2
x20[31] i_instruction[15] net46[31] net47[31] net42 net45[31] mux2
x20[30] i_instruction[15] net46[30] net47[30] net42 net45[30] mux2
x20[29] i_instruction[15] net46[29] net47[29] net42 net45[29] mux2
x20[28] i_instruction[15] net46[28] net47[28] net42 net45[28] mux2
x20[27] i_instruction[15] net46[27] net47[27] net42 net45[27] mux2
x20[26] i_instruction[15] net46[26] net47[26] net42 net45[26] mux2
x20[25] i_instruction[15] net46[25] net47[25] net42 net45[25] mux2
x20[24] i_instruction[15] net46[24] net47[24] net42 net45[24] mux2
x20[23] i_instruction[15] net46[23] net47[23] net42 net45[23] mux2
x20[22] i_instruction[15] net46[22] net47[22] net42 net45[22] mux2
x20[21] i_instruction[15] net46[21] net47[21] net42 net45[21] mux2
x20[20] i_instruction[15] net46[20] net47[20] net42 net45[20] mux2
x20[19] i_instruction[15] net46[19] net47[19] net42 net45[19] mux2
x20[18] i_instruction[15] net46[18] net47[18] net42 net45[18] mux2
x20[17] i_instruction[15] net46[17] net47[17] net42 net45[17] mux2
x20[16] i_instruction[15] net46[16] net47[16] net42 net45[16] mux2
x20[15] i_instruction[15] net46[15] net47[15] net42 net45[15] mux2
x20[14] i_instruction[15] net46[14] net47[14] net42 net45[14] mux2
x20[13] i_instruction[15] net46[13] net47[13] net42 net45[13] mux2
x20[12] i_instruction[15] net46[12] net47[12] net42 net45[12] mux2
x20[11] i_instruction[15] net46[11] net47[11] net42 net45[11] mux2
x20[10] i_instruction[15] net46[10] net47[10] net42 net45[10] mux2
x20[9] i_instruction[15] net46[9] net47[9] net42 net45[9] mux2
x20[8] i_instruction[15] net46[8] net47[8] net42 net45[8] mux2
x20[7] i_instruction[15] net46[7] net47[7] net42 net45[7] mux2
x20[6] i_instruction[15] net46[6] net47[6] net42 net45[6] mux2
x20[5] i_instruction[15] net46[5] net47[5] net42 net45[5] mux2
x20[4] i_instruction[15] net46[4] net47[4] net42 net45[4] mux2
x20[3] i_instruction[15] net46[3] net47[3] net42 net45[3] mux2
x20[2] i_instruction[15] net46[2] net47[2] net42 net45[2] mux2
x20[1] i_instruction[15] net46[1] net47[1] net42 net45[1] mux2
x20[0] i_instruction[15] net46[0] net47[0] net42 net45[0] mux2
x31 i_instruction[15] VSS VSS VCC VCC net42 sky130_fd_sc_hd__inv_1
x21[32] i_instruction[14] VSS net45[32] net43 VSS mux2
x21[31] i_instruction[14] VSS net45[31] net43 VSS mux2
x21[30] i_instruction[14] VSS net45[30] net43 VSS mux2
x21[29] i_instruction[14] VSS net45[29] net43 VSS mux2
x21[28] i_instruction[14] VSS net45[28] net43 VSS mux2
x21[27] i_instruction[14] i_instruction[3] net45[27] net43 VSS mux2
x21[26] i_instruction[14] i_instruction[2] net45[26] net43 VSS mux2
x21[25] i_instruction[14] i_instruction[12] net45[25] net43 VSS mux2
x21[24] i_instruction[14] i_instruction[6] net45[24] net43 i_instruction[6] mux2
x21[23] i_instruction[14] i_instruction[5] net45[23] net43 i_instruction[5] mux2
x21[22] i_instruction[14] i_instruction[4] net45[22] net43 i_instruction[4] mux2
x21[21] i_instruction[14] VSS net45[21] net43 i_instruction[3] mux2
x21[20] i_instruction[14] VSS net45[20] net43 i_instruction[2] mux2
x21[19] i_instruction[14] VSS net45[19] net43 i_instruction[11] mux2
x21[18] i_instruction[14] VSS net45[18] net43 i_instruction[10] mux2
x21[17] i_instruction[14] VSS net45[17] net43 i_instruction[9] mux2
x21[16] i_instruction[14] VCC net45[16] net43 i_instruction[8] mux2
x21[15] i_instruction[14] VSS net45[15] net43 i_instruction[7] mux2
x21[14] i_instruction[14] VSS net45[14] net43 VSS mux2
x21[13] i_instruction[14] VCC net45[13] net43 VSS mux2
x21[12] i_instruction[14] VSS net45[12] net43 VCC mux2
x21[11] i_instruction[14] i_instruction[11] net45[11] net43 i_instruction[11] mux2
x21[10] i_instruction[14] i_instruction[10] net45[10] net43 i_instruction[10] mux2
x21[9] i_instruction[14] i_instruction[9] net45[9] net43 i_instruction[9] mux2
x21[8] i_instruction[14] i_instruction[8] net45[8] net43 i_instruction[8] mux2
x21[7] i_instruction[14] i_instruction[7] net45[7] net43 i_instruction[7] mux2
x21[6] i_instruction[14] VSS net45[6] net43 VSS mux2
x21[5] i_instruction[14] VSS net45[5] net43 VSS mux2
x21[4] i_instruction[14] VSS net45[4] net43 VCC mux2
x21[3] i_instruction[14] VSS net45[3] net43 VSS mux2
x21[2] i_instruction[14] VSS net45[2] net43 VSS mux2
x21[1] i_instruction[14] VCC net45[1] net43 VCC mux2
x21[0] i_instruction[14] VCC net45[0] net43 VCC mux2
x32 i_instruction[14] VSS VSS VCC VCC net43 sky130_fd_sc_hd__inv_1
x22[32] i_instruction[14] VSS net46[32] net44 net50[32] mux2
x22[31] i_instruction[14] VSS net46[31] net44 net50[31] mux2
x22[30] i_instruction[14] VSS net46[30] net44 net50[30] mux2
x22[29] i_instruction[14] VSS net46[29] net44 net50[29] mux2
x22[28] i_instruction[14] VSS net46[28] net44 net50[28] mux2
x22[27] i_instruction[14] i_instruction[8] net46[27] net44 net50[27] mux2
x22[26] i_instruction[14] i_instruction[7] net46[26] net44 net50[26] mux2
x22[25] i_instruction[14] i_instruction[12] net46[25] net44 net50[25] mux2
x22[24] i_instruction[14] i_instruction[6] net46[24] net44 net50[24] mux2
x22[23] i_instruction[14] i_instruction[5] net46[23] net44 net50[23] mux2
x22[22] i_instruction[14] i_instruction[4] net46[22] net44 net50[22] mux2
x22[21] i_instruction[14] i_instruction[3] net46[21] net44 net50[21] mux2
x22[20] i_instruction[14] i_instruction[2] net46[20] net44 net50[20] mux2
x22[19] i_instruction[14] VSS net46[19] net44 net50[19] mux2
x22[18] i_instruction[14] VSS net46[18] net44 net50[18] mux2
x22[17] i_instruction[14] VSS net46[17] net44 net50[17] mux2
x22[16] i_instruction[14] VCC net46[16] net44 net50[16] mux2
x22[15] i_instruction[14] VSS net46[15] net44 net50[15] mux2
x22[14] i_instruction[14] VSS net46[14] net44 net50[14] mux2
x22[13] i_instruction[14] VCC net46[13] net44 net50[13] mux2
x22[12] i_instruction[14] VSS net46[12] net44 net50[12] mux2
x22[11] i_instruction[14] i_instruction[11] net46[11] net44 net50[11] mux2
x22[10] i_instruction[14] i_instruction[10] net46[10] net44 net50[10] mux2
x22[9] i_instruction[14] i_instruction[9] net46[9] net44 net50[9] mux2
x22[8] i_instruction[14] VSS net46[8] net44 net50[8] mux2
x22[7] i_instruction[14] VSS net46[7] net44 net50[7] mux2
x22[6] i_instruction[14] VSS net46[6] net44 net50[6] mux2
x22[5] i_instruction[14] VCC net46[5] net44 net50[5] mux2
x22[4] i_instruction[14] VSS net46[4] net44 net50[4] mux2
x22[3] i_instruction[14] VSS net46[3] net44 net50[3] mux2
x22[2] i_instruction[14] VSS net46[2] net44 net50[2] mux2
x22[1] i_instruction[14] VCC net46[1] net44 net50[1] mux2
x22[0] i_instruction[14] VCC net46[0] net44 net50[0] mux2
x33 i_instruction[14] VSS VSS VCC VCC net44 sky130_fd_sc_hd__inv_1
x23[32] i_instruction[12] net56[32] net50[32] net49 net54[32] mux2
x23[31] i_instruction[12] net56[31] net50[31] net49 net54[31] mux2
x23[30] i_instruction[12] net56[30] net50[30] net49 net54[30] mux2
x23[29] i_instruction[12] net56[29] net50[29] net49 net54[29] mux2
x23[28] i_instruction[12] net56[28] net50[28] net49 net54[28] mux2
x23[27] i_instruction[12] net56[27] net50[27] net49 net54[27] mux2
x23[26] i_instruction[12] net56[26] net50[26] net49 net54[26] mux2
x23[25] i_instruction[12] net56[25] net50[25] net49 net54[25] mux2
x23[24] i_instruction[12] net56[24] net50[24] net49 net54[24] mux2
x23[23] i_instruction[12] net56[23] net50[23] net49 net54[23] mux2
x23[22] i_instruction[12] net56[22] net50[22] net49 net54[22] mux2
x23[21] i_instruction[12] net56[21] net50[21] net49 net54[21] mux2
x23[20] i_instruction[12] net56[20] net50[20] net49 net54[20] mux2
x23[19] i_instruction[12] net56[19] net50[19] net49 net54[19] mux2
x23[18] i_instruction[12] net56[18] net50[18] net49 net54[18] mux2
x23[17] i_instruction[12] net56[17] net50[17] net49 net54[17] mux2
x23[16] i_instruction[12] net56[16] net50[16] net49 net54[16] mux2
x23[15] i_instruction[12] net56[15] net50[15] net49 net54[15] mux2
x23[14] i_instruction[12] net56[14] net50[14] net49 net54[14] mux2
x23[13] i_instruction[12] net56[13] net50[13] net49 net54[13] mux2
x23[12] i_instruction[12] net56[12] net50[12] net49 net54[12] mux2
x23[11] i_instruction[12] net56[11] net50[11] net49 net54[11] mux2
x23[10] i_instruction[12] net56[10] net50[10] net49 net54[10] mux2
x23[9] i_instruction[12] net56[9] net50[9] net49 net54[9] mux2
x23[8] i_instruction[12] net56[8] net50[8] net49 net54[8] mux2
x23[7] i_instruction[12] net56[7] net50[7] net49 net54[7] mux2
x23[6] i_instruction[12] net56[6] net50[6] net49 net54[6] mux2
x23[5] i_instruction[12] net56[5] net50[5] net49 net54[5] mux2
x23[4] i_instruction[12] net56[4] net50[4] net49 net54[4] mux2
x23[3] i_instruction[12] net56[3] net50[3] net49 net54[3] mux2
x23[2] i_instruction[12] net56[2] net50[2] net49 net54[2] mux2
x23[1] i_instruction[12] net56[1] net50[1] net49 net54[1] mux2
x23[0] i_instruction[12] net56[0] net50[0] net49 net54[0] mux2
x34 i_instruction[12] VSS VSS VCC VCC net49 sky130_fd_sc_hd__inv_1
x24[32] net51 VSS net54[32] net52 VSS mux2
x24[31] net51 VSS net54[31] net52 VSS mux2
x24[30] net51 VSS net54[30] net52 VSS mux2
x24[29] net51 VSS net54[29] net52 VSS mux2
x24[28] net51 VSS net54[28] net52 VSS mux2
x24[27] net51 VSS net54[27] net52 VSS mux2
x24[26] net51 VSS net54[26] net52 VSS mux2
x24[25] net51 VSS net54[25] net52 VSS mux2
x24[24] net51 i_instruction[6] net54[24] net52 VSS mux2
x24[23] net51 i_instruction[5] net54[23] net52 VSS mux2
x24[22] net51 i_instruction[4] net54[22] net52 VSS mux2
x24[21] net51 i_instruction[3] net54[21] net52 VSS mux2
x24[20] net51 i_instruction[2] net54[20] net52 VSS mux2
x24[19] net51 VSS net54[19] net52 i_instruction[11] mux2
x24[18] net51 VSS net54[18] net52 i_instruction[10] mux2
x24[17] net51 VSS net54[17] net52 i_instruction[9] mux2
x24[16] net51 VSS net54[16] net52 i_instruction[8] mux2
x24[15] net51 VSS net54[15] net52 i_instruction[7] mux2
x24[14] net51 VSS net54[14] net52 VSS mux2
x24[13] net51 VSS net54[13] net52 VSS mux2
x24[12] net51 VSS net54[12] net52 VSS mux2
x24[11] net51 i_instruction[11] net54[11] net52 VSS mux2
x24[10] net51 i_instruction[10] net54[10] net52 VSS mux2
x24[9] net51 i_instruction[9] net54[9] net52 VSS mux2
x24[8] net51 i_instruction[8] net54[8] net52 VSS mux2
x24[7] net51 i_instruction[7] net54[7] net52 VSS mux2
x24[6] net51 VSS net54[6] net52 VCC mux2
x24[5] net51 VCC net54[5] net52 VCC mux2
x24[4] net51 VCC net54[4] net52 VSS mux2
x24[3] net51 VSS net54[3] net52 VSS mux2
x24[2] net51 VSS net54[2] net52 VCC mux2
x24[1] net51 VCC net54[1] net52 VCC mux2
x24[0] net51 VCC net54[0] net52 VCC mux2
x35 net51 VSS VSS VCC VCC net52 sky130_fd_sc_hd__inv_1
x36 i_instruction[6] i_instruction[5] i_instruction[4] VSS VSS VCC VCC net67 sky130_fd_sc_hd__or3_1
x37 i_instruction[3] i_instruction[2] VSS VSS VCC VCC net53 sky130_fd_sc_hd__or2_1
x38 net67 net53 VSS VSS VCC VCC net51 sky130_fd_sc_hd__or2_1
x25[32] net51 VSS net56[32] net55 net59[32] mux2
x25[31] net51 VSS net56[31] net55 net59[31] mux2
x25[30] net51 VSS net56[30] net55 net59[30] mux2
x25[29] net51 VSS net56[29] net55 net59[29] mux2
x25[28] net51 VSS net56[28] net55 net59[28] mux2
x25[27] net51 VSS net56[27] net55 net59[27] mux2
x25[26] net51 VSS net56[26] net55 net59[26] mux2
x25[25] net51 VSS net56[25] net55 net59[25] mux2
x25[24] net51 i_instruction[6] net56[24] net55 net59[24] mux2
x25[23] net51 i_instruction[5] net56[23] net55 net59[23] mux2
x25[22] net51 i_instruction[4] net56[22] net55 net59[22] mux2
x25[21] net51 i_instruction[3] net56[21] net55 net59[21] mux2
x25[20] net51 i_instruction[2] net56[20] net55 net59[20] mux2
x25[19] net51 i_instruction[11] net56[19] net55 net59[19] mux2
x25[18] net51 i_instruction[10] net56[18] net55 net59[18] mux2
x25[17] net51 i_instruction[9] net56[17] net55 net59[17] mux2
x25[16] net51 i_instruction[8] net56[16] net55 net59[16] mux2
x25[15] net51 i_instruction[7] net56[15] net55 net59[15] mux2
x25[14] net51 VSS net56[14] net55 net59[14] mux2
x25[13] net51 VSS net56[13] net55 net59[13] mux2
x25[12] net51 VSS net56[12] net55 net59[12] mux2
x25[11] net51 i_instruction[11] net56[11] net55 net59[11] mux2
x25[10] net51 i_instruction[10] net56[10] net55 net59[10] mux2
x25[9] net51 i_instruction[9] net56[9] net55 net59[9] mux2
x25[8] net51 i_instruction[8] net56[8] net55 net59[8] mux2
x25[7] net51 i_instruction[7] net56[7] net55 net59[7] mux2
x25[6] net51 VSS net56[6] net55 net59[6] mux2
x25[5] net51 VCC net56[5] net55 net59[5] mux2
x25[4] net51 VCC net56[4] net55 net59[4] mux2
x25[3] net51 VSS net56[3] net55 net59[3] mux2
x25[2] net51 VSS net56[2] net55 net59[2] mux2
x25[1] net51 VCC net56[1] net55 net59[1] mux2
x25[0] net51 VCC net56[0] net55 net59[0] mux2
x39 net51 VSS VSS VCC VCC net55 sky130_fd_sc_hd__inv_1
x26[32] net57 VSS net59[32] net58 VSS mux2
x26[31] net57 VSS net59[31] net58 VSS mux2
x26[30] net57 VSS net59[30] net58 VSS mux2
x26[29] net57 VSS net59[29] net58 VSS mux2
x26[28] net57 VSS net59[28] net58 VSS mux2
x26[27] net57 VSS net59[27] net58 VSS mux2
x26[26] net57 VSS net59[26] net58 VSS mux2
x26[25] net57 VSS net59[25] net58 VSS mux2
x26[24] net57 VSS net59[24] net58 VSS mux2
x26[23] net57 VSS net59[23] net58 VSS mux2
x26[22] net57 VSS net59[22] net58 VSS mux2
x26[21] net57 VSS net59[21] net58 VSS mux2
x26[20] net57 VCC net59[20] net58 VSS mux2
x26[19] net57 VSS net59[19] net58 i_instruction[11] mux2
x26[18] net57 VSS net59[18] net58 i_instruction[10] mux2
x26[17] net57 VSS net59[17] net58 i_instruction[9] mux2
x26[16] net57 VSS net59[16] net58 i_instruction[8] mux2
x26[15] net57 VSS net59[15] net58 i_instruction[7] mux2
x26[14] net57 VSS net59[14] net58 VSS mux2
x26[13] net57 VSS net59[13] net58 VSS mux2
x26[12] net57 VSS net59[12] net58 VSS mux2
x26[11] net57 VSS net59[11] net58 VSS mux2
x26[10] net57 VSS net59[10] net58 VSS mux2
x26[9] net57 VSS net59[9] net58 VSS mux2
x26[8] net57 VSS net59[8] net58 VSS mux2
x26[7] net57 VSS net59[7] net58 VCC mux2
x26[6] net57 VCC net59[6] net58 VCC mux2
x26[5] net57 VCC net59[5] net58 VCC mux2
x26[4] net57 VCC net59[4] net58 VSS mux2
x26[3] net57 VSS net59[3] net58 VSS mux2
x26[2] net57 VSS net59[2] net58 VCC mux2
x26[1] net57 VCC net59[1] net58 VCC mux2
x26[0] net57 VCC net59[0] net58 VCC mux2
x40 net57 VSS VSS VCC VCC net58 sky130_fd_sc_hd__inv_1
x41 i_instruction[11] i_instruction[10] i_instruction[9] VSS VSS VCC VCC net68
+ sky130_fd_sc_hd__or3_1
x42 i_instruction[8] i_instruction[7] VSS VSS VCC VCC net60 sky130_fd_sc_hd__or2_1
x43 net68 net60 VSS VSS VCC VCC net57 sky130_fd_sc_hd__nor2_1
**.ends

* expanding   symbol:  ../../elements/logic/mux2.sym # of pins=5
** sym_path: /media/FlexRV32/asic/elements/logic/mux2.sym
** sch_path: /media/FlexRV32/asic/elements/logic/mux2.sch
.subckt mux2 s0 d0 Y s1 d1
*.ipin s0
*.ipin d0
*.ipin s1
*.ipin d1
*.opin Y
x1 s0 d0 VSS VSS VCC VCC net1 sky130_fd_sc_hd__nand2_1
x2 s1 d1 VSS VSS VCC VCC net2 sky130_fd_sc_hd__nand2_1
x3 net1 net2 VSS VSS VCC VCC Y sky130_fd_sc_hd__nand2_1
.ends

.GLOBAL VSS
.GLOBAL VCC
.end
