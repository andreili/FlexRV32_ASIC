* ROM data
* Generated file, don't change!
* Selection buffer
xSELBUF0 SEL VSS VSS VCC VCC SEL0 sky130_fd_sc_hd__inv_1
xSELBUF1 SEL0 VSS VSS VCC VCC SEL1 sky130_fd_sc_hd__inv_2
xSELBUF2 SEL1 VSS VSS VCC VCC SEL2 sky130_fd_sc_hd__inv_8
* Bitlines pull-up
XPM[0] BL[0] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[1] BL[1] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[2] BL[2] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[3] BL[3] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[4] BL[4] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[5] BL[5] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[6] BL[6] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[7] BL[7] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[8] BL[8] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[9] BL[9] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[10] BL[10] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[11] BL[11] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[12] BL[12] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[13] BL[13] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[14] BL[14] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[15] BL[15] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[16] BL[16] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[17] BL[17] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[18] BL[18] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[19] BL[19] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[20] BL[20] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[21] BL[21] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[22] BL[22] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[23] BL[23] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[24] BL[24] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[25] BL[25] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[26] BL[26] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[27] BL[27] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[28] BL[28] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[29] BL[29] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[30] BL[30] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[31] BL[31] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[32] BL[32] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[33] BL[33] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[34] BL[34] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[35] BL[35] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[36] BL[36] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[37] BL[37] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[38] BL[38] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[39] BL[39] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[40] BL[40] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[41] BL[41] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[42] BL[42] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[43] BL[43] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[44] BL[44] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[45] BL[45] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[46] BL[46] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[47] BL[47] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[48] BL[48] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[49] BL[49] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[50] BL[50] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[51] BL[51] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[52] BL[52] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[53] BL[53] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[54] BL[54] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[55] BL[55] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[56] BL[56] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[57] BL[57] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[58] BL[58] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[59] BL[59] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[60] BL[60] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[61] BL[61] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[62] BL[62] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[63] BL[63] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[64] BL[64] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[65] BL[65] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[66] BL[66] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[67] BL[67] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[68] BL[68] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[69] BL[69] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[70] BL[70] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[71] BL[71] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[72] BL[72] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[73] BL[73] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[74] BL[74] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[75] BL[75] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[76] BL[76] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[77] BL[77] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[78] BL[78] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[79] BL[79] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[80] BL[80] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[81] BL[81] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[82] BL[82] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[83] BL[83] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[84] BL[84] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[85] BL[85] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[86] BL[86] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[87] BL[87] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[88] BL[88] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[89] BL[89] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[90] BL[90] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[91] BL[91] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[92] BL[92] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[93] BL[93] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[94] BL[94] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[95] BL[95] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[96] BL[96] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[97] BL[97] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[98] BL[98] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[99] BL[99] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[100] BL[100] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[101] BL[101] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[102] BL[102] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[103] BL[103] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[104] BL[104] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[105] BL[105] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[106] BL[106] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[107] BL[107] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[108] BL[108] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[109] BL[109] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[110] BL[110] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[111] BL[111] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[112] BL[112] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[113] BL[113] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[114] BL[114] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[115] BL[115] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[116] BL[116] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[117] BL[117] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[118] BL[118] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[119] BL[119] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[120] BL[120] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[121] BL[121] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[122] BL[122] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[123] BL[123] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[124] BL[124] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[125] BL[125] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[126] BL[126] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
XPM[127] BL[127] SEL2 VCC VCC sky130_fd_pr__pfet_01v8_hvt w=650000u l=150000u
* Word lines buffers
xBUF0_0[0] ROW[0] VSS VSS VCC VCC WL0[0] sky130_fd_sc_hd__inv_2
xBUF0_0[1] ROW[1] VSS VSS VCC VCC WL0[1] sky130_fd_sc_hd__inv_2
xBUF0_0[2] ROW[2] VSS VSS VCC VCC WL0[2] sky130_fd_sc_hd__inv_2
xBUF0_0[3] ROW[3] VSS VSS VCC VCC WL0[3] sky130_fd_sc_hd__inv_2
xBUF0_0[4] ROW[4] VSS VSS VCC VCC WL0[4] sky130_fd_sc_hd__inv_2
xBUF0_0[5] ROW[5] VSS VSS VCC VCC WL0[5] sky130_fd_sc_hd__inv_2
xBUF0_0[6] ROW[6] VSS VSS VCC VCC WL0[6] sky130_fd_sc_hd__inv_2
xBUF0_0[7] ROW[7] VSS VSS VCC VCC WL0[7] sky130_fd_sc_hd__inv_2
xBUF0_0[8] ROW[8] VSS VSS VCC VCC WL0[8] sky130_fd_sc_hd__inv_2
xBUF0_0[9] ROW[9] VSS VSS VCC VCC WL0[9] sky130_fd_sc_hd__inv_2
xBUF0_0[10] ROW[10] VSS VSS VCC VCC WL0[10] sky130_fd_sc_hd__inv_2
xBUF0_0[11] ROW[11] VSS VSS VCC VCC WL0[11] sky130_fd_sc_hd__inv_2
xBUF0_0[12] ROW[12] VSS VSS VCC VCC WL0[12] sky130_fd_sc_hd__inv_2
xBUF0_0[13] ROW[13] VSS VSS VCC VCC WL0[13] sky130_fd_sc_hd__inv_2
xBUF0_0[14] ROW[14] VSS VSS VCC VCC WL0[14] sky130_fd_sc_hd__inv_2
xBUF0_0[15] ROW[15] VSS VSS VCC VCC WL0[15] sky130_fd_sc_hd__inv_2
xBUF0_0[16] ROW[16] VSS VSS VCC VCC WL0[16] sky130_fd_sc_hd__inv_2
xBUF0_0[17] ROW[17] VSS VSS VCC VCC WL0[17] sky130_fd_sc_hd__inv_2
xBUF0_0[18] ROW[18] VSS VSS VCC VCC WL0[18] sky130_fd_sc_hd__inv_2
xBUF0_0[19] ROW[19] VSS VSS VCC VCC WL0[19] sky130_fd_sc_hd__inv_2
xBUF0_0[20] ROW[20] VSS VSS VCC VCC WL0[20] sky130_fd_sc_hd__inv_2
xBUF0_0[21] ROW[21] VSS VSS VCC VCC WL0[21] sky130_fd_sc_hd__inv_2
xBUF0_0[22] ROW[22] VSS VSS VCC VCC WL0[22] sky130_fd_sc_hd__inv_2
xBUF0_0[23] ROW[23] VSS VSS VCC VCC WL0[23] sky130_fd_sc_hd__inv_2
xBUF0_0[24] ROW[24] VSS VSS VCC VCC WL0[24] sky130_fd_sc_hd__inv_2
xBUF0_0[25] ROW[25] VSS VSS VCC VCC WL0[25] sky130_fd_sc_hd__inv_2
xBUF0_0[26] ROW[26] VSS VSS VCC VCC WL0[26] sky130_fd_sc_hd__inv_2
xBUF0_0[27] ROW[27] VSS VSS VCC VCC WL0[27] sky130_fd_sc_hd__inv_2
xBUF0_0[28] ROW[28] VSS VSS VCC VCC WL0[28] sky130_fd_sc_hd__inv_2
xBUF0_0[29] ROW[29] VSS VSS VCC VCC WL0[29] sky130_fd_sc_hd__inv_2
xBUF0_0[30] ROW[30] VSS VSS VCC VCC WL0[30] sky130_fd_sc_hd__inv_2
xBUF0_0[31] ROW[31] VSS VSS VCC VCC WL0[31] sky130_fd_sc_hd__inv_2
xBUF0_0[32] ROW[32] VSS VSS VCC VCC WL0[32] sky130_fd_sc_hd__inv_2
xBUF0_0[33] ROW[33] VSS VSS VCC VCC WL0[33] sky130_fd_sc_hd__inv_2
xBUF0_0[34] ROW[34] VSS VSS VCC VCC WL0[34] sky130_fd_sc_hd__inv_2
xBUF0_0[35] ROW[35] VSS VSS VCC VCC WL0[35] sky130_fd_sc_hd__inv_2
xBUF0_0[36] ROW[36] VSS VSS VCC VCC WL0[36] sky130_fd_sc_hd__inv_2
xBUF0_0[37] ROW[37] VSS VSS VCC VCC WL0[37] sky130_fd_sc_hd__inv_2
xBUF0_0[38] ROW[38] VSS VSS VCC VCC WL0[38] sky130_fd_sc_hd__inv_2
xBUF0_0[39] ROW[39] VSS VSS VCC VCC WL0[39] sky130_fd_sc_hd__inv_2
xBUF0_0[40] ROW[40] VSS VSS VCC VCC WL0[40] sky130_fd_sc_hd__inv_2
xBUF0_0[41] ROW[41] VSS VSS VCC VCC WL0[41] sky130_fd_sc_hd__inv_2
xBUF0_0[42] ROW[42] VSS VSS VCC VCC WL0[42] sky130_fd_sc_hd__inv_2
xBUF0_0[43] ROW[43] VSS VSS VCC VCC WL0[43] sky130_fd_sc_hd__inv_2
xBUF0_0[44] ROW[44] VSS VSS VCC VCC WL0[44] sky130_fd_sc_hd__inv_2
xBUF0_0[45] ROW[45] VSS VSS VCC VCC WL0[45] sky130_fd_sc_hd__inv_2
xBUF0_0[46] ROW[46] VSS VSS VCC VCC WL0[46] sky130_fd_sc_hd__inv_2
xBUF0_0[47] ROW[47] VSS VSS VCC VCC WL0[47] sky130_fd_sc_hd__inv_2
xBUF0_0[48] ROW[48] VSS VSS VCC VCC WL0[48] sky130_fd_sc_hd__inv_2
xBUF0_0[49] ROW[49] VSS VSS VCC VCC WL0[49] sky130_fd_sc_hd__inv_2
xBUF0_0[50] ROW[50] VSS VSS VCC VCC WL0[50] sky130_fd_sc_hd__inv_2
xBUF0_0[51] ROW[51] VSS VSS VCC VCC WL0[51] sky130_fd_sc_hd__inv_2
xBUF0_0[52] ROW[52] VSS VSS VCC VCC WL0[52] sky130_fd_sc_hd__inv_2
xBUF0_0[53] ROW[53] VSS VSS VCC VCC WL0[53] sky130_fd_sc_hd__inv_2
xBUF0_0[54] ROW[54] VSS VSS VCC VCC WL0[54] sky130_fd_sc_hd__inv_2
xBUF0_0[55] ROW[55] VSS VSS VCC VCC WL0[55] sky130_fd_sc_hd__inv_2
xBUF0_0[56] ROW[56] VSS VSS VCC VCC WL0[56] sky130_fd_sc_hd__inv_2
xBUF0_0[57] ROW[57] VSS VSS VCC VCC WL0[57] sky130_fd_sc_hd__inv_2
xBUF0_0[58] ROW[58] VSS VSS VCC VCC WL0[58] sky130_fd_sc_hd__inv_2
xBUF0_0[59] ROW[59] VSS VSS VCC VCC WL0[59] sky130_fd_sc_hd__inv_2
xBUF0_0[60] ROW[60] VSS VSS VCC VCC WL0[60] sky130_fd_sc_hd__inv_2
xBUF0_0[61] ROW[61] VSS VSS VCC VCC WL0[61] sky130_fd_sc_hd__inv_2
xBUF0_0[62] ROW[62] VSS VSS VCC VCC WL0[62] sky130_fd_sc_hd__inv_2
xBUF0_0[63] ROW[63] VSS VSS VCC VCC WL0[63] sky130_fd_sc_hd__inv_2
xBUF0_0[64] ROW[64] VSS VSS VCC VCC WL0[64] sky130_fd_sc_hd__inv_2
xBUF0_0[65] ROW[65] VSS VSS VCC VCC WL0[65] sky130_fd_sc_hd__inv_2
xBUF0_0[66] ROW[66] VSS VSS VCC VCC WL0[66] sky130_fd_sc_hd__inv_2
xBUF0_0[67] ROW[67] VSS VSS VCC VCC WL0[67] sky130_fd_sc_hd__inv_2
xBUF0_0[68] ROW[68] VSS VSS VCC VCC WL0[68] sky130_fd_sc_hd__inv_2
xBUF0_0[69] ROW[69] VSS VSS VCC VCC WL0[69] sky130_fd_sc_hd__inv_2
xBUF0_0[70] ROW[70] VSS VSS VCC VCC WL0[70] sky130_fd_sc_hd__inv_2
xBUF0_0[71] ROW[71] VSS VSS VCC VCC WL0[71] sky130_fd_sc_hd__inv_2
xBUF0_0[72] ROW[72] VSS VSS VCC VCC WL0[72] sky130_fd_sc_hd__inv_2
xBUF0_0[73] ROW[73] VSS VSS VCC VCC WL0[73] sky130_fd_sc_hd__inv_2
xBUF0_0[74] ROW[74] VSS VSS VCC VCC WL0[74] sky130_fd_sc_hd__inv_2
xBUF0_0[75] ROW[75] VSS VSS VCC VCC WL0[75] sky130_fd_sc_hd__inv_2
xBUF0_0[76] ROW[76] VSS VSS VCC VCC WL0[76] sky130_fd_sc_hd__inv_2
xBUF0_0[77] ROW[77] VSS VSS VCC VCC WL0[77] sky130_fd_sc_hd__inv_2
xBUF0_0[78] ROW[78] VSS VSS VCC VCC WL0[78] sky130_fd_sc_hd__inv_2
xBUF0_0[79] ROW[79] VSS VSS VCC VCC WL0[79] sky130_fd_sc_hd__inv_2
xBUF0_0[80] ROW[80] VSS VSS VCC VCC WL0[80] sky130_fd_sc_hd__inv_2
xBUF0_0[81] ROW[81] VSS VSS VCC VCC WL0[81] sky130_fd_sc_hd__inv_2
xBUF0_0[82] ROW[82] VSS VSS VCC VCC WL0[82] sky130_fd_sc_hd__inv_2
xBUF0_0[83] ROW[83] VSS VSS VCC VCC WL0[83] sky130_fd_sc_hd__inv_2
xBUF0_0[84] ROW[84] VSS VSS VCC VCC WL0[84] sky130_fd_sc_hd__inv_2
xBUF0_0[85] ROW[85] VSS VSS VCC VCC WL0[85] sky130_fd_sc_hd__inv_2
xBUF0_0[86] ROW[86] VSS VSS VCC VCC WL0[86] sky130_fd_sc_hd__inv_2
xBUF0_0[87] ROW[87] VSS VSS VCC VCC WL0[87] sky130_fd_sc_hd__inv_2
xBUF0_0[88] ROW[88] VSS VSS VCC VCC WL0[88] sky130_fd_sc_hd__inv_2
xBUF0_0[89] ROW[89] VSS VSS VCC VCC WL0[89] sky130_fd_sc_hd__inv_2
xBUF0_0[90] ROW[90] VSS VSS VCC VCC WL0[90] sky130_fd_sc_hd__inv_2
xBUF0_0[91] ROW[91] VSS VSS VCC VCC WL0[91] sky130_fd_sc_hd__inv_2
xBUF0_0[92] ROW[92] VSS VSS VCC VCC WL0[92] sky130_fd_sc_hd__inv_2
xBUF0_0[93] ROW[93] VSS VSS VCC VCC WL0[93] sky130_fd_sc_hd__inv_2
xBUF0_0[94] ROW[94] VSS VSS VCC VCC WL0[94] sky130_fd_sc_hd__inv_2
xBUF0_0[95] ROW[95] VSS VSS VCC VCC WL0[95] sky130_fd_sc_hd__inv_2
xBUF0_0[96] ROW[96] VSS VSS VCC VCC WL0[96] sky130_fd_sc_hd__inv_2
xBUF0_0[97] ROW[97] VSS VSS VCC VCC WL0[97] sky130_fd_sc_hd__inv_2
xBUF0_0[98] ROW[98] VSS VSS VCC VCC WL0[98] sky130_fd_sc_hd__inv_2
xBUF0_0[99] ROW[99] VSS VSS VCC VCC WL0[99] sky130_fd_sc_hd__inv_2
xBUF0_0[100] ROW[100] VSS VSS VCC VCC WL0[100] sky130_fd_sc_hd__inv_2
xBUF0_0[101] ROW[101] VSS VSS VCC VCC WL0[101] sky130_fd_sc_hd__inv_2
xBUF0_0[102] ROW[102] VSS VSS VCC VCC WL0[102] sky130_fd_sc_hd__inv_2
xBUF0_0[103] ROW[103] VSS VSS VCC VCC WL0[103] sky130_fd_sc_hd__inv_2
xBUF0_0[104] ROW[104] VSS VSS VCC VCC WL0[104] sky130_fd_sc_hd__inv_2
xBUF0_0[105] ROW[105] VSS VSS VCC VCC WL0[105] sky130_fd_sc_hd__inv_2
xBUF0_0[106] ROW[106] VSS VSS VCC VCC WL0[106] sky130_fd_sc_hd__inv_2
xBUF0_0[107] ROW[107] VSS VSS VCC VCC WL0[107] sky130_fd_sc_hd__inv_2
xBUF0_0[108] ROW[108] VSS VSS VCC VCC WL0[108] sky130_fd_sc_hd__inv_2
xBUF0_0[109] ROW[109] VSS VSS VCC VCC WL0[109] sky130_fd_sc_hd__inv_2
xBUF0_0[110] ROW[110] VSS VSS VCC VCC WL0[110] sky130_fd_sc_hd__inv_2
xBUF0_0[111] ROW[111] VSS VSS VCC VCC WL0[111] sky130_fd_sc_hd__inv_2
xBUF0_0[112] ROW[112] VSS VSS VCC VCC WL0[112] sky130_fd_sc_hd__inv_2
xBUF0_0[113] ROW[113] VSS VSS VCC VCC WL0[113] sky130_fd_sc_hd__inv_2
xBUF0_0[114] ROW[114] VSS VSS VCC VCC WL0[114] sky130_fd_sc_hd__inv_2
xBUF0_0[115] ROW[115] VSS VSS VCC VCC WL0[115] sky130_fd_sc_hd__inv_2
xBUF0_0[116] ROW[116] VSS VSS VCC VCC WL0[116] sky130_fd_sc_hd__inv_2
xBUF0_0[117] ROW[117] VSS VSS VCC VCC WL0[117] sky130_fd_sc_hd__inv_2
xBUF0_0[118] ROW[118] VSS VSS VCC VCC WL0[118] sky130_fd_sc_hd__inv_2
xBUF0_0[119] ROW[119] VSS VSS VCC VCC WL0[119] sky130_fd_sc_hd__inv_2
xBUF0_0[120] ROW[120] VSS VSS VCC VCC WL0[120] sky130_fd_sc_hd__inv_2
xBUF0_0[121] ROW[121] VSS VSS VCC VCC WL0[121] sky130_fd_sc_hd__inv_2
xBUF0_0[122] ROW[122] VSS VSS VCC VCC WL0[122] sky130_fd_sc_hd__inv_2
xBUF0_0[123] ROW[123] VSS VSS VCC VCC WL0[123] sky130_fd_sc_hd__inv_2
xBUF0_0[124] ROW[124] VSS VSS VCC VCC WL0[124] sky130_fd_sc_hd__inv_2
xBUF0_0[125] ROW[125] VSS VSS VCC VCC WL0[125] sky130_fd_sc_hd__inv_2
xBUF0_0[126] ROW[126] VSS VSS VCC VCC WL0[126] sky130_fd_sc_hd__inv_2
xBUF0_0[127] ROW[127] VSS VSS VCC VCC WL0[127] sky130_fd_sc_hd__inv_2
xBUF0_0[128] ROW[128] VSS VSS VCC VCC WL0[128] sky130_fd_sc_hd__inv_2
xBUF0_0[129] ROW[129] VSS VSS VCC VCC WL0[129] sky130_fd_sc_hd__inv_2
xBUF0_0[130] ROW[130] VSS VSS VCC VCC WL0[130] sky130_fd_sc_hd__inv_2
xBUF0_0[131] ROW[131] VSS VSS VCC VCC WL0[131] sky130_fd_sc_hd__inv_2
xBUF0_0[132] ROW[132] VSS VSS VCC VCC WL0[132] sky130_fd_sc_hd__inv_2
xBUF0_0[133] ROW[133] VSS VSS VCC VCC WL0[133] sky130_fd_sc_hd__inv_2
xBUF0_0[134] ROW[134] VSS VSS VCC VCC WL0[134] sky130_fd_sc_hd__inv_2
xBUF0_0[135] ROW[135] VSS VSS VCC VCC WL0[135] sky130_fd_sc_hd__inv_2
xBUF0_0[136] ROW[136] VSS VSS VCC VCC WL0[136] sky130_fd_sc_hd__inv_2
xBUF0_0[137] ROW[137] VSS VSS VCC VCC WL0[137] sky130_fd_sc_hd__inv_2
xBUF0_0[138] ROW[138] VSS VSS VCC VCC WL0[138] sky130_fd_sc_hd__inv_2
xBUF0_0[139] ROW[139] VSS VSS VCC VCC WL0[139] sky130_fd_sc_hd__inv_2
xBUF0_0[140] ROW[140] VSS VSS VCC VCC WL0[140] sky130_fd_sc_hd__inv_2
xBUF0_0[141] ROW[141] VSS VSS VCC VCC WL0[141] sky130_fd_sc_hd__inv_2
xBUF0_0[142] ROW[142] VSS VSS VCC VCC WL0[142] sky130_fd_sc_hd__inv_2
xBUF0_0[143] ROW[143] VSS VSS VCC VCC WL0[143] sky130_fd_sc_hd__inv_2
xBUF0_0[144] ROW[144] VSS VSS VCC VCC WL0[144] sky130_fd_sc_hd__inv_2
xBUF0_0[145] ROW[145] VSS VSS VCC VCC WL0[145] sky130_fd_sc_hd__inv_2
xBUF0_0[146] ROW[146] VSS VSS VCC VCC WL0[146] sky130_fd_sc_hd__inv_2
xBUF0_0[147] ROW[147] VSS VSS VCC VCC WL0[147] sky130_fd_sc_hd__inv_2
xBUF0_0[148] ROW[148] VSS VSS VCC VCC WL0[148] sky130_fd_sc_hd__inv_2
xBUF0_0[149] ROW[149] VSS VSS VCC VCC WL0[149] sky130_fd_sc_hd__inv_2
xBUF0_0[150] ROW[150] VSS VSS VCC VCC WL0[150] sky130_fd_sc_hd__inv_2
xBUF0_0[151] ROW[151] VSS VSS VCC VCC WL0[151] sky130_fd_sc_hd__inv_2
xBUF0_0[152] ROW[152] VSS VSS VCC VCC WL0[152] sky130_fd_sc_hd__inv_2
xBUF0_0[153] ROW[153] VSS VSS VCC VCC WL0[153] sky130_fd_sc_hd__inv_2
xBUF0_0[154] ROW[154] VSS VSS VCC VCC WL0[154] sky130_fd_sc_hd__inv_2
xBUF0_0[155] ROW[155] VSS VSS VCC VCC WL0[155] sky130_fd_sc_hd__inv_2
xBUF0_0[156] ROW[156] VSS VSS VCC VCC WL0[156] sky130_fd_sc_hd__inv_2
xBUF0_0[157] ROW[157] VSS VSS VCC VCC WL0[157] sky130_fd_sc_hd__inv_2
xBUF0_0[158] ROW[158] VSS VSS VCC VCC WL0[158] sky130_fd_sc_hd__inv_2
xBUF0_0[159] ROW[159] VSS VSS VCC VCC WL0[159] sky130_fd_sc_hd__inv_2
xBUF0_0[160] ROW[160] VSS VSS VCC VCC WL0[160] sky130_fd_sc_hd__inv_2
xBUF0_0[161] ROW[161] VSS VSS VCC VCC WL0[161] sky130_fd_sc_hd__inv_2
xBUF0_0[162] ROW[162] VSS VSS VCC VCC WL0[162] sky130_fd_sc_hd__inv_2
xBUF0_0[163] ROW[163] VSS VSS VCC VCC WL0[163] sky130_fd_sc_hd__inv_2
xBUF0_0[164] ROW[164] VSS VSS VCC VCC WL0[164] sky130_fd_sc_hd__inv_2
xBUF0_0[165] ROW[165] VSS VSS VCC VCC WL0[165] sky130_fd_sc_hd__inv_2
xBUF0_0[166] ROW[166] VSS VSS VCC VCC WL0[166] sky130_fd_sc_hd__inv_2
xBUF0_0[167] ROW[167] VSS VSS VCC VCC WL0[167] sky130_fd_sc_hd__inv_2
xBUF0_0[168] ROW[168] VSS VSS VCC VCC WL0[168] sky130_fd_sc_hd__inv_2
xBUF0_0[169] ROW[169] VSS VSS VCC VCC WL0[169] sky130_fd_sc_hd__inv_2
xBUF0_0[170] ROW[170] VSS VSS VCC VCC WL0[170] sky130_fd_sc_hd__inv_2
xBUF0_0[171] ROW[171] VSS VSS VCC VCC WL0[171] sky130_fd_sc_hd__inv_2
xBUF0_0[172] ROW[172] VSS VSS VCC VCC WL0[172] sky130_fd_sc_hd__inv_2
xBUF0_0[173] ROW[173] VSS VSS VCC VCC WL0[173] sky130_fd_sc_hd__inv_2
xBUF0_0[174] ROW[174] VSS VSS VCC VCC WL0[174] sky130_fd_sc_hd__inv_2
xBUF0_0[175] ROW[175] VSS VSS VCC VCC WL0[175] sky130_fd_sc_hd__inv_2
xBUF0_0[176] ROW[176] VSS VSS VCC VCC WL0[176] sky130_fd_sc_hd__inv_2
xBUF0_0[177] ROW[177] VSS VSS VCC VCC WL0[177] sky130_fd_sc_hd__inv_2
xBUF0_0[178] ROW[178] VSS VSS VCC VCC WL0[178] sky130_fd_sc_hd__inv_2
xBUF0_0[179] ROW[179] VSS VSS VCC VCC WL0[179] sky130_fd_sc_hd__inv_2
xBUF0_0[180] ROW[180] VSS VSS VCC VCC WL0[180] sky130_fd_sc_hd__inv_2
xBUF0_0[181] ROW[181] VSS VSS VCC VCC WL0[181] sky130_fd_sc_hd__inv_2
xBUF0_0[182] ROW[182] VSS VSS VCC VCC WL0[182] sky130_fd_sc_hd__inv_2
xBUF0_0[183] ROW[183] VSS VSS VCC VCC WL0[183] sky130_fd_sc_hd__inv_2
xBUF0_0[184] ROW[184] VSS VSS VCC VCC WL0[184] sky130_fd_sc_hd__inv_2
xBUF0_0[185] ROW[185] VSS VSS VCC VCC WL0[185] sky130_fd_sc_hd__inv_2
xBUF0_0[186] ROW[186] VSS VSS VCC VCC WL0[186] sky130_fd_sc_hd__inv_2
xBUF0_0[187] ROW[187] VSS VSS VCC VCC WL0[187] sky130_fd_sc_hd__inv_2
xBUF0_0[188] ROW[188] VSS VSS VCC VCC WL0[188] sky130_fd_sc_hd__inv_2
xBUF0_0[189] ROW[189] VSS VSS VCC VCC WL0[189] sky130_fd_sc_hd__inv_2
xBUF0_0[190] ROW[190] VSS VSS VCC VCC WL0[190] sky130_fd_sc_hd__inv_2
xBUF0_0[191] ROW[191] VSS VSS VCC VCC WL0[191] sky130_fd_sc_hd__inv_2
xBUF0_0[192] ROW[192] VSS VSS VCC VCC WL0[192] sky130_fd_sc_hd__inv_2
xBUF0_0[193] ROW[193] VSS VSS VCC VCC WL0[193] sky130_fd_sc_hd__inv_2
xBUF0_0[194] ROW[194] VSS VSS VCC VCC WL0[194] sky130_fd_sc_hd__inv_2
xBUF0_0[195] ROW[195] VSS VSS VCC VCC WL0[195] sky130_fd_sc_hd__inv_2
xBUF0_0[196] ROW[196] VSS VSS VCC VCC WL0[196] sky130_fd_sc_hd__inv_2
xBUF0_0[197] ROW[197] VSS VSS VCC VCC WL0[197] sky130_fd_sc_hd__inv_2
xBUF0_0[198] ROW[198] VSS VSS VCC VCC WL0[198] sky130_fd_sc_hd__inv_2
xBUF0_0[199] ROW[199] VSS VSS VCC VCC WL0[199] sky130_fd_sc_hd__inv_2
xBUF0_0[200] ROW[200] VSS VSS VCC VCC WL0[200] sky130_fd_sc_hd__inv_2
xBUF0_0[201] ROW[201] VSS VSS VCC VCC WL0[201] sky130_fd_sc_hd__inv_2
xBUF0_0[202] ROW[202] VSS VSS VCC VCC WL0[202] sky130_fd_sc_hd__inv_2
xBUF0_0[203] ROW[203] VSS VSS VCC VCC WL0[203] sky130_fd_sc_hd__inv_2
xBUF0_0[204] ROW[204] VSS VSS VCC VCC WL0[204] sky130_fd_sc_hd__inv_2
xBUF0_0[205] ROW[205] VSS VSS VCC VCC WL0[205] sky130_fd_sc_hd__inv_2
xBUF0_0[206] ROW[206] VSS VSS VCC VCC WL0[206] sky130_fd_sc_hd__inv_2
xBUF0_0[207] ROW[207] VSS VSS VCC VCC WL0[207] sky130_fd_sc_hd__inv_2
xBUF0_0[208] ROW[208] VSS VSS VCC VCC WL0[208] sky130_fd_sc_hd__inv_2
xBUF0_0[209] ROW[209] VSS VSS VCC VCC WL0[209] sky130_fd_sc_hd__inv_2
xBUF0_0[210] ROW[210] VSS VSS VCC VCC WL0[210] sky130_fd_sc_hd__inv_2
xBUF0_0[211] ROW[211] VSS VSS VCC VCC WL0[211] sky130_fd_sc_hd__inv_2
xBUF0_0[212] ROW[212] VSS VSS VCC VCC WL0[212] sky130_fd_sc_hd__inv_2
xBUF0_0[213] ROW[213] VSS VSS VCC VCC WL0[213] sky130_fd_sc_hd__inv_2
xBUF0_0[214] ROW[214] VSS VSS VCC VCC WL0[214] sky130_fd_sc_hd__inv_2
xBUF0_0[215] ROW[215] VSS VSS VCC VCC WL0[215] sky130_fd_sc_hd__inv_2
xBUF0_0[216] ROW[216] VSS VSS VCC VCC WL0[216] sky130_fd_sc_hd__inv_2
xBUF0_0[217] ROW[217] VSS VSS VCC VCC WL0[217] sky130_fd_sc_hd__inv_2
xBUF0_0[218] ROW[218] VSS VSS VCC VCC WL0[218] sky130_fd_sc_hd__inv_2
xBUF0_0[219] ROW[219] VSS VSS VCC VCC WL0[219] sky130_fd_sc_hd__inv_2
xBUF0_0[220] ROW[220] VSS VSS VCC VCC WL0[220] sky130_fd_sc_hd__inv_2
xBUF0_0[221] ROW[221] VSS VSS VCC VCC WL0[221] sky130_fd_sc_hd__inv_2
xBUF0_0[222] ROW[222] VSS VSS VCC VCC WL0[222] sky130_fd_sc_hd__inv_2
xBUF0_0[223] ROW[223] VSS VSS VCC VCC WL0[223] sky130_fd_sc_hd__inv_2
xBUF0_0[224] ROW[224] VSS VSS VCC VCC WL0[224] sky130_fd_sc_hd__inv_2
xBUF0_0[225] ROW[225] VSS VSS VCC VCC WL0[225] sky130_fd_sc_hd__inv_2
xBUF0_0[226] ROW[226] VSS VSS VCC VCC WL0[226] sky130_fd_sc_hd__inv_2
xBUF0_0[227] ROW[227] VSS VSS VCC VCC WL0[227] sky130_fd_sc_hd__inv_2
xBUF0_0[228] ROW[228] VSS VSS VCC VCC WL0[228] sky130_fd_sc_hd__inv_2
xBUF0_0[229] ROW[229] VSS VSS VCC VCC WL0[229] sky130_fd_sc_hd__inv_2
xBUF0_0[230] ROW[230] VSS VSS VCC VCC WL0[230] sky130_fd_sc_hd__inv_2
xBUF0_0[231] ROW[231] VSS VSS VCC VCC WL0[231] sky130_fd_sc_hd__inv_2
xBUF0_0[232] ROW[232] VSS VSS VCC VCC WL0[232] sky130_fd_sc_hd__inv_2
xBUF0_0[233] ROW[233] VSS VSS VCC VCC WL0[233] sky130_fd_sc_hd__inv_2
xBUF0_0[234] ROW[234] VSS VSS VCC VCC WL0[234] sky130_fd_sc_hd__inv_2
xBUF0_0[235] ROW[235] VSS VSS VCC VCC WL0[235] sky130_fd_sc_hd__inv_2
xBUF0_0[236] ROW[236] VSS VSS VCC VCC WL0[236] sky130_fd_sc_hd__inv_2
xBUF0_0[237] ROW[237] VSS VSS VCC VCC WL0[237] sky130_fd_sc_hd__inv_2
xBUF0_0[238] ROW[238] VSS VSS VCC VCC WL0[238] sky130_fd_sc_hd__inv_2
xBUF0_0[239] ROW[239] VSS VSS VCC VCC WL0[239] sky130_fd_sc_hd__inv_2
xBUF0_0[240] ROW[240] VSS VSS VCC VCC WL0[240] sky130_fd_sc_hd__inv_2
xBUF0_0[241] ROW[241] VSS VSS VCC VCC WL0[241] sky130_fd_sc_hd__inv_2
xBUF0_0[242] ROW[242] VSS VSS VCC VCC WL0[242] sky130_fd_sc_hd__inv_2
xBUF0_0[243] ROW[243] VSS VSS VCC VCC WL0[243] sky130_fd_sc_hd__inv_2
xBUF0_0[244] ROW[244] VSS VSS VCC VCC WL0[244] sky130_fd_sc_hd__inv_2
xBUF0_0[245] ROW[245] VSS VSS VCC VCC WL0[245] sky130_fd_sc_hd__inv_2
xBUF0_0[246] ROW[246] VSS VSS VCC VCC WL0[246] sky130_fd_sc_hd__inv_2
xBUF0_0[247] ROW[247] VSS VSS VCC VCC WL0[247] sky130_fd_sc_hd__inv_2
xBUF0_0[248] ROW[248] VSS VSS VCC VCC WL0[248] sky130_fd_sc_hd__inv_2
xBUF0_0[249] ROW[249] VSS VSS VCC VCC WL0[249] sky130_fd_sc_hd__inv_2
xBUF0_0[250] ROW[250] VSS VSS VCC VCC WL0[250] sky130_fd_sc_hd__inv_2
xBUF0_0[251] ROW[251] VSS VSS VCC VCC WL0[251] sky130_fd_sc_hd__inv_2
xBUF0_0[252] ROW[252] VSS VSS VCC VCC WL0[252] sky130_fd_sc_hd__inv_2
xBUF0_0[253] ROW[253] VSS VSS VCC VCC WL0[253] sky130_fd_sc_hd__inv_2
xBUF0_0[254] ROW[254] VSS VSS VCC VCC WL0[254] sky130_fd_sc_hd__inv_2
xBUF0_0[255] ROW[255] VSS VSS VCC VCC WL0[255] sky130_fd_sc_hd__inv_2
* Column driver buffers
xCBUF0[0] COL[0] VSS VSS VCC VCC COL_B0_n[0] sky130_fd_sc_hd__inv_1
xCBUF0p0[0] COL_B0_n[0] VSS VSS VCC VCC COL_B10_p[0] sky130_fd_sc_hd__inv_1
xCBUF0n0[0] COL_B10_p[0] VSS VSS VCC VCC COL_B10_n[0] sky130_fd_sc_hd__inv_1
xCBUF0p1[0] COL_B0_n[0] VSS VSS VCC VCC COL_B11_p[0] sky130_fd_sc_hd__inv_1
xCBUF0n1[0] COL_B11_p[0] VSS VSS VCC VCC COL_B11_n[0] sky130_fd_sc_hd__inv_1
xCBUF0p2[0] COL_B0_n[0] VSS VSS VCC VCC COL_B12_p[0] sky130_fd_sc_hd__inv_1
xCBUF0n2[0] COL_B12_p[0] VSS VSS VCC VCC COL_B12_n[0] sky130_fd_sc_hd__inv_1
xCBUF0p3[0] COL_B0_n[0] VSS VSS VCC VCC COL_B13_p[0] sky130_fd_sc_hd__inv_1
xCBUF0n3[0] COL_B13_p[0] VSS VSS VCC VCC COL_B13_n[0] sky130_fd_sc_hd__inv_1
xCBUF0[1] COL[1] VSS VSS VCC VCC COL_B0_n[1] sky130_fd_sc_hd__inv_1
xCBUF0p0[1] COL_B0_n[1] VSS VSS VCC VCC COL_B10_p[1] sky130_fd_sc_hd__inv_1
xCBUF0n0[1] COL_B10_p[1] VSS VSS VCC VCC COL_B10_n[1] sky130_fd_sc_hd__inv_1
xCBUF0p1[1] COL_B0_n[1] VSS VSS VCC VCC COL_B11_p[1] sky130_fd_sc_hd__inv_1
xCBUF0n1[1] COL_B11_p[1] VSS VSS VCC VCC COL_B11_n[1] sky130_fd_sc_hd__inv_1
xCBUF0p2[1] COL_B0_n[1] VSS VSS VCC VCC COL_B12_p[1] sky130_fd_sc_hd__inv_1
xCBUF0n2[1] COL_B12_p[1] VSS VSS VCC VCC COL_B12_n[1] sky130_fd_sc_hd__inv_1
xCBUF0p3[1] COL_B0_n[1] VSS VSS VCC VCC COL_B13_p[1] sky130_fd_sc_hd__inv_1
xCBUF0n3[1] COL_B13_p[1] VSS VSS VCC VCC COL_B13_n[1] sky130_fd_sc_hd__inv_1
xCBUF0[2] COL[2] VSS VSS VCC VCC COL_B0_n[2] sky130_fd_sc_hd__inv_1
xCBUF0p0[2] COL_B0_n[2] VSS VSS VCC VCC COL_B10_p[2] sky130_fd_sc_hd__inv_1
xCBUF0n0[2] COL_B10_p[2] VSS VSS VCC VCC COL_B10_n[2] sky130_fd_sc_hd__inv_1
xCBUF0p1[2] COL_B0_n[2] VSS VSS VCC VCC COL_B11_p[2] sky130_fd_sc_hd__inv_1
xCBUF0n1[2] COL_B11_p[2] VSS VSS VCC VCC COL_B11_n[2] sky130_fd_sc_hd__inv_1
xCBUF0p2[2] COL_B0_n[2] VSS VSS VCC VCC COL_B12_p[2] sky130_fd_sc_hd__inv_1
xCBUF0n2[2] COL_B12_p[2] VSS VSS VCC VCC COL_B12_n[2] sky130_fd_sc_hd__inv_1
xCBUF0p3[2] COL_B0_n[2] VSS VSS VCC VCC COL_B13_p[2] sky130_fd_sc_hd__inv_1
xCBUF0n3[2] COL_B13_p[2] VSS VSS VCC VCC COL_B13_n[2] sky130_fd_sc_hd__inv_1
xCBUF0[3] COL[3] VSS VSS VCC VCC COL_B0_n[3] sky130_fd_sc_hd__inv_1
xCBUF0p0[3] COL_B0_n[3] VSS VSS VCC VCC COL_B10_p[3] sky130_fd_sc_hd__inv_1
xCBUF0n0[3] COL_B10_p[3] VSS VSS VCC VCC COL_B10_n[3] sky130_fd_sc_hd__inv_1
xCBUF0p1[3] COL_B0_n[3] VSS VSS VCC VCC COL_B11_p[3] sky130_fd_sc_hd__inv_1
xCBUF0n1[3] COL_B11_p[3] VSS VSS VCC VCC COL_B11_n[3] sky130_fd_sc_hd__inv_1
xCBUF0p2[3] COL_B0_n[3] VSS VSS VCC VCC COL_B12_p[3] sky130_fd_sc_hd__inv_1
xCBUF0n2[3] COL_B12_p[3] VSS VSS VCC VCC COL_B12_n[3] sky130_fd_sc_hd__inv_1
xCBUF0p3[3] COL_B0_n[3] VSS VSS VCC VCC COL_B13_p[3] sky130_fd_sc_hd__inv_1
xCBUF0n3[3] COL_B13_p[3] VSS VSS VCC VCC COL_B13_n[3] sky130_fd_sc_hd__inv_1
* Data array
* addr: 0x0
XM1 VSS WL0[0] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2 VSS WL0[0] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3 VSS WL0[0] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4 VSS WL0[0] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5 VSS WL0[0] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6 VSS WL0[0] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7 VSS WL0[0] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8 VSS WL0[0] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM9 VSS WL0[0] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM10 VSS WL0[0] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM11 VSS WL0[0] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM12 VSS WL0[0] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM13 VSS WL0[0] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM14 VSS WL0[0] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM15 VSS WL0[0] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM16 VSS WL0[0] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM17 VSS WL0[0] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM18 VSS WL0[0] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM19 VSS WL0[0] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM20 VSS WL0[0] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM21 VSS WL0[0] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM22 VSS WL0[0] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM23 VSS WL0[0] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM24 VSS WL0[0] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM25 VSS WL0[0] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM26 VSS WL0[0] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM27 VSS WL0[0] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM28 VSS WL0[0] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM29 VSS WL0[0] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM30 VSS WL0[0] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM31 VSS WL0[0] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM32 VSS WL0[0] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM33 VSS WL0[0] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM34 VSS WL0[0] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM35 VSS WL0[0] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM36 VSS WL0[0] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM37 VSS WL0[0] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x10
XM38 VSS WL0[1] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM39 VSS WL0[1] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM40 VSS WL0[1] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM41 VSS WL0[1] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM42 VSS WL0[1] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM43 VSS WL0[1] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM44 VSS WL0[1] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM45 VSS WL0[1] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM46 VSS WL0[1] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM47 VSS WL0[1] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM48 VSS WL0[1] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM49 VSS WL0[1] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM50 VSS WL0[1] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM51 VSS WL0[1] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM52 VSS WL0[1] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM53 VSS WL0[1] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM54 VSS WL0[1] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM55 VSS WL0[1] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM56 VSS WL0[1] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM57 VSS WL0[1] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM58 VSS WL0[1] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM59 VSS WL0[1] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM60 VSS WL0[1] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM61 VSS WL0[1] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM62 VSS WL0[1] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM63 VSS WL0[1] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM64 VSS WL0[1] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM65 VSS WL0[1] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM66 VSS WL0[1] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM67 VSS WL0[1] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM68 VSS WL0[1] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM69 VSS WL0[1] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM70 VSS WL0[1] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM71 VSS WL0[1] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM72 VSS WL0[1] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM73 VSS WL0[1] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM74 VSS WL0[1] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM75 VSS WL0[1] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM76 VSS WL0[1] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x20
XM77 VSS WL0[2] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM78 VSS WL0[2] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM79 VSS WL0[2] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM80 VSS WL0[2] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM81 VSS WL0[2] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM82 VSS WL0[2] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM83 VSS WL0[2] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM84 VSS WL0[2] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM85 VSS WL0[2] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM86 VSS WL0[2] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM87 VSS WL0[2] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM88 VSS WL0[2] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM89 VSS WL0[2] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM90 VSS WL0[2] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM91 VSS WL0[2] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM92 VSS WL0[2] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM93 VSS WL0[2] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM94 VSS WL0[2] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM95 VSS WL0[2] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM96 VSS WL0[2] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM97 VSS WL0[2] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM98 VSS WL0[2] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM99 VSS WL0[2] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM100 VSS WL0[2] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM101 VSS WL0[2] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM102 VSS WL0[2] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM103 VSS WL0[2] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM104 VSS WL0[2] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM105 VSS WL0[2] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM106 VSS WL0[2] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM107 VSS WL0[2] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM108 VSS WL0[2] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM109 VSS WL0[2] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM110 VSS WL0[2] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM111 VSS WL0[2] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM112 VSS WL0[2] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM113 VSS WL0[2] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM114 VSS WL0[2] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM115 VSS WL0[2] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM116 VSS WL0[2] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM117 VSS WL0[2] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM118 VSS WL0[2] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM119 VSS WL0[2] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM120 VSS WL0[2] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM121 VSS WL0[2] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM122 VSS WL0[2] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM123 VSS WL0[2] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x30
XM124 VSS WL0[3] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM125 VSS WL0[3] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM126 VSS WL0[3] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM127 VSS WL0[3] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM128 VSS WL0[3] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM129 VSS WL0[3] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM130 VSS WL0[3] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM131 VSS WL0[3] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM132 VSS WL0[3] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM133 VSS WL0[3] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM134 VSS WL0[3] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM135 VSS WL0[3] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM136 VSS WL0[3] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM137 VSS WL0[3] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM138 VSS WL0[3] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM139 VSS WL0[3] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM140 VSS WL0[3] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM141 VSS WL0[3] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM142 VSS WL0[3] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM143 VSS WL0[3] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM144 VSS WL0[3] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM145 VSS WL0[3] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM146 VSS WL0[3] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM147 VSS WL0[3] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM148 VSS WL0[3] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM149 VSS WL0[3] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM150 VSS WL0[3] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM151 VSS WL0[3] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM152 VSS WL0[3] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM153 VSS WL0[3] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM154 VSS WL0[3] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM155 VSS WL0[3] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM156 VSS WL0[3] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM157 VSS WL0[3] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM158 VSS WL0[3] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM159 VSS WL0[3] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM160 VSS WL0[3] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM161 VSS WL0[3] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM162 VSS WL0[3] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM163 VSS WL0[3] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM164 VSS WL0[3] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM165 VSS WL0[3] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM166 VSS WL0[3] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM167 VSS WL0[3] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM168 VSS WL0[3] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM169 VSS WL0[3] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM170 VSS WL0[3] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM171 VSS WL0[3] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x40
XM172 VSS WL0[4] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM173 VSS WL0[4] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM174 VSS WL0[4] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM175 VSS WL0[4] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM176 VSS WL0[4] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM177 VSS WL0[4] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM178 VSS WL0[4] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM179 VSS WL0[4] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM180 VSS WL0[4] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM181 VSS WL0[4] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM182 VSS WL0[4] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM183 VSS WL0[4] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM184 VSS WL0[4] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM185 VSS WL0[4] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM186 VSS WL0[4] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM187 VSS WL0[4] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM188 VSS WL0[4] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM189 VSS WL0[4] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM190 VSS WL0[4] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM191 VSS WL0[4] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM192 VSS WL0[4] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM193 VSS WL0[4] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM194 VSS WL0[4] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM195 VSS WL0[4] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM196 VSS WL0[4] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM197 VSS WL0[4] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM198 VSS WL0[4] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM199 VSS WL0[4] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM200 VSS WL0[4] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM201 VSS WL0[4] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM202 VSS WL0[4] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM203 VSS WL0[4] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM204 VSS WL0[4] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM205 VSS WL0[4] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM206 VSS WL0[4] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM207 VSS WL0[4] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM208 VSS WL0[4] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM209 VSS WL0[4] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM210 VSS WL0[4] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x50
XM211 VSS WL0[5] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM212 VSS WL0[5] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM213 VSS WL0[5] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM214 VSS WL0[5] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM215 VSS WL0[5] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM216 VSS WL0[5] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM217 VSS WL0[5] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM218 VSS WL0[5] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM219 VSS WL0[5] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM220 VSS WL0[5] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM221 VSS WL0[5] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM222 VSS WL0[5] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM223 VSS WL0[5] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM224 VSS WL0[5] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM225 VSS WL0[5] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM226 VSS WL0[5] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM227 VSS WL0[5] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM228 VSS WL0[5] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM229 VSS WL0[5] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM230 VSS WL0[5] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM231 VSS WL0[5] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM232 VSS WL0[5] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM233 VSS WL0[5] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM234 VSS WL0[5] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM235 VSS WL0[5] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM236 VSS WL0[5] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM237 VSS WL0[5] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM238 VSS WL0[5] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM239 VSS WL0[5] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM240 VSS WL0[5] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM241 VSS WL0[5] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM242 VSS WL0[5] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM243 VSS WL0[5] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM244 VSS WL0[5] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM245 VSS WL0[5] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM246 VSS WL0[5] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM247 VSS WL0[5] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM248 VSS WL0[5] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM249 VSS WL0[5] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM250 VSS WL0[5] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM251 VSS WL0[5] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM252 VSS WL0[5] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM253 VSS WL0[5] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM254 VSS WL0[5] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM255 VSS WL0[5] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM256 VSS WL0[5] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM257 VSS WL0[5] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM258 VSS WL0[5] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x60
XM259 VSS WL0[6] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM260 VSS WL0[6] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM261 VSS WL0[6] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM262 VSS WL0[6] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM263 VSS WL0[6] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM264 VSS WL0[6] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM265 VSS WL0[6] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM266 VSS WL0[6] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM267 VSS WL0[6] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM268 VSS WL0[6] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM269 VSS WL0[6] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM270 VSS WL0[6] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM271 VSS WL0[6] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM272 VSS WL0[6] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM273 VSS WL0[6] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM274 VSS WL0[6] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM275 VSS WL0[6] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM276 VSS WL0[6] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM277 VSS WL0[6] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM278 VSS WL0[6] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM279 VSS WL0[6] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM280 VSS WL0[6] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM281 VSS WL0[6] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM282 VSS WL0[6] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM283 VSS WL0[6] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM284 VSS WL0[6] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM285 VSS WL0[6] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM286 VSS WL0[6] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM287 VSS WL0[6] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM288 VSS WL0[6] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM289 VSS WL0[6] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM290 VSS WL0[6] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM291 VSS WL0[6] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM292 VSS WL0[6] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM293 VSS WL0[6] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM294 VSS WL0[6] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM295 VSS WL0[6] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM296 VSS WL0[6] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM297 VSS WL0[6] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM298 VSS WL0[6] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM299 VSS WL0[6] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM300 VSS WL0[6] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM301 VSS WL0[6] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM302 VSS WL0[6] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM303 VSS WL0[6] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM304 VSS WL0[6] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM305 VSS WL0[6] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM306 VSS WL0[6] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM307 VSS WL0[6] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM308 VSS WL0[6] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM309 VSS WL0[6] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM310 VSS WL0[6] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM311 VSS WL0[6] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM312 VSS WL0[6] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM313 VSS WL0[6] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x70
XM314 VSS WL0[7] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM315 VSS WL0[7] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM316 VSS WL0[7] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM317 VSS WL0[7] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM318 VSS WL0[7] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM319 VSS WL0[7] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM320 VSS WL0[7] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM321 VSS WL0[7] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM322 VSS WL0[7] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM323 VSS WL0[7] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM324 VSS WL0[7] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM325 VSS WL0[7] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM326 VSS WL0[7] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM327 VSS WL0[7] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM328 VSS WL0[7] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM329 VSS WL0[7] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM330 VSS WL0[7] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM331 VSS WL0[7] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM332 VSS WL0[7] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM333 VSS WL0[7] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM334 VSS WL0[7] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM335 VSS WL0[7] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM336 VSS WL0[7] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM337 VSS WL0[7] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM338 VSS WL0[7] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM339 VSS WL0[7] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM340 VSS WL0[7] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM341 VSS WL0[7] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM342 VSS WL0[7] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM343 VSS WL0[7] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM344 VSS WL0[7] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM345 VSS WL0[7] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM346 VSS WL0[7] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM347 VSS WL0[7] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM348 VSS WL0[7] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM349 VSS WL0[7] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM350 VSS WL0[7] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM351 VSS WL0[7] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM352 VSS WL0[7] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM353 VSS WL0[7] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM354 VSS WL0[7] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM355 VSS WL0[7] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM356 VSS WL0[7] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM357 VSS WL0[7] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM358 VSS WL0[7] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM359 VSS WL0[7] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x80
XM360 VSS WL0[8] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM361 VSS WL0[8] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM362 VSS WL0[8] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM363 VSS WL0[8] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM364 VSS WL0[8] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM365 VSS WL0[8] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM366 VSS WL0[8] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM367 VSS WL0[8] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM368 VSS WL0[8] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM369 VSS WL0[8] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM370 VSS WL0[8] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM371 VSS WL0[8] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM372 VSS WL0[8] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM373 VSS WL0[8] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM374 VSS WL0[8] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM375 VSS WL0[8] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM376 VSS WL0[8] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM377 VSS WL0[8] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM378 VSS WL0[8] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM379 VSS WL0[8] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM380 VSS WL0[8] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM381 VSS WL0[8] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM382 VSS WL0[8] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM383 VSS WL0[8] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM384 VSS WL0[8] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM385 VSS WL0[8] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM386 VSS WL0[8] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM387 VSS WL0[8] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM388 VSS WL0[8] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM389 VSS WL0[8] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM390 VSS WL0[8] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM391 VSS WL0[8] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM392 VSS WL0[8] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM393 VSS WL0[8] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM394 VSS WL0[8] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM395 VSS WL0[8] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM396 VSS WL0[8] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM397 VSS WL0[8] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM398 VSS WL0[8] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM399 VSS WL0[8] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM400 VSS WL0[8] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM401 VSS WL0[8] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM402 VSS WL0[8] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM403 VSS WL0[8] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM404 VSS WL0[8] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x90
XM405 VSS WL0[9] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM406 VSS WL0[9] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM407 VSS WL0[9] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM408 VSS WL0[9] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM409 VSS WL0[9] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM410 VSS WL0[9] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM411 VSS WL0[9] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM412 VSS WL0[9] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM413 VSS WL0[9] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM414 VSS WL0[9] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM415 VSS WL0[9] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM416 VSS WL0[9] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM417 VSS WL0[9] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM418 VSS WL0[9] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM419 VSS WL0[9] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM420 VSS WL0[9] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM421 VSS WL0[9] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM422 VSS WL0[9] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM423 VSS WL0[9] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM424 VSS WL0[9] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM425 VSS WL0[9] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM426 VSS WL0[9] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM427 VSS WL0[9] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM428 VSS WL0[9] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM429 VSS WL0[9] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM430 VSS WL0[9] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM431 VSS WL0[9] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM432 VSS WL0[9] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM433 VSS WL0[9] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM434 VSS WL0[9] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM435 VSS WL0[9] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM436 VSS WL0[9] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM437 VSS WL0[9] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM438 VSS WL0[9] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM439 VSS WL0[9] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM440 VSS WL0[9] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM441 VSS WL0[9] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM442 VSS WL0[9] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM443 VSS WL0[9] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM444 VSS WL0[9] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM445 VSS WL0[9] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM446 VSS WL0[9] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM447 VSS WL0[9] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM448 VSS WL0[9] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM449 VSS WL0[9] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM450 VSS WL0[9] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM451 VSS WL0[9] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM452 VSS WL0[9] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM453 VSS WL0[9] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM454 VSS WL0[9] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM455 VSS WL0[9] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM456 VSS WL0[9] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM457 VSS WL0[9] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM458 VSS WL0[9] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM459 VSS WL0[9] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM460 VSS WL0[9] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM461 VSS WL0[9] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM462 VSS WL0[9] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM463 VSS WL0[9] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM464 VSS WL0[9] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM465 VSS WL0[9] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM466 VSS WL0[9] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM467 VSS WL0[9] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0xa0
XM468 VSS WL0[10] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM469 VSS WL0[10] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM470 VSS WL0[10] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM471 VSS WL0[10] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM472 VSS WL0[10] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM473 VSS WL0[10] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM474 VSS WL0[10] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM475 VSS WL0[10] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM476 VSS WL0[10] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM477 VSS WL0[10] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM478 VSS WL0[10] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM479 VSS WL0[10] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM480 VSS WL0[10] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM481 VSS WL0[10] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM482 VSS WL0[10] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM483 VSS WL0[10] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM484 VSS WL0[10] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM485 VSS WL0[10] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM486 VSS WL0[10] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM487 VSS WL0[10] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM488 VSS WL0[10] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM489 VSS WL0[10] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM490 VSS WL0[10] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM491 VSS WL0[10] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM492 VSS WL0[10] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM493 VSS WL0[10] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM494 VSS WL0[10] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM495 VSS WL0[10] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM496 VSS WL0[10] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM497 VSS WL0[10] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM498 VSS WL0[10] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM499 VSS WL0[10] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM500 VSS WL0[10] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM501 VSS WL0[10] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM502 VSS WL0[10] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM503 VSS WL0[10] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM504 VSS WL0[10] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM505 VSS WL0[10] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM506 VSS WL0[10] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM507 VSS WL0[10] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM508 VSS WL0[10] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM509 VSS WL0[10] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM510 VSS WL0[10] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM511 VSS WL0[10] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM512 VSS WL0[10] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM513 VSS WL0[10] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM514 VSS WL0[10] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM515 VSS WL0[10] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM516 VSS WL0[10] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM517 VSS WL0[10] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM518 VSS WL0[10] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM519 VSS WL0[10] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM520 VSS WL0[10] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM521 VSS WL0[10] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM522 VSS WL0[10] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM523 VSS WL0[10] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM524 VSS WL0[10] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM525 VSS WL0[10] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM526 VSS WL0[10] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM527 VSS WL0[10] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM528 VSS WL0[10] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM529 VSS WL0[10] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM530 VSS WL0[10] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM531 VSS WL0[10] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM532 VSS WL0[10] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM533 VSS WL0[10] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0xb0
XM534 VSS WL0[11] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM535 VSS WL0[11] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM536 VSS WL0[11] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM537 VSS WL0[11] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM538 VSS WL0[11] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM539 VSS WL0[11] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM540 VSS WL0[11] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM541 VSS WL0[11] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM542 VSS WL0[11] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM543 VSS WL0[11] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM544 VSS WL0[11] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM545 VSS WL0[11] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM546 VSS WL0[11] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM547 VSS WL0[11] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM548 VSS WL0[11] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM549 VSS WL0[11] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM550 VSS WL0[11] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM551 VSS WL0[11] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM552 VSS WL0[11] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM553 VSS WL0[11] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM554 VSS WL0[11] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM555 VSS WL0[11] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM556 VSS WL0[11] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM557 VSS WL0[11] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM558 VSS WL0[11] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM559 VSS WL0[11] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM560 VSS WL0[11] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM561 VSS WL0[11] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM562 VSS WL0[11] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM563 VSS WL0[11] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM564 VSS WL0[11] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM565 VSS WL0[11] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM566 VSS WL0[11] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM567 VSS WL0[11] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM568 VSS WL0[11] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM569 VSS WL0[11] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM570 VSS WL0[11] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM571 VSS WL0[11] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM572 VSS WL0[11] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM573 VSS WL0[11] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM574 VSS WL0[11] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM575 VSS WL0[11] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM576 VSS WL0[11] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0xc0
XM577 VSS WL0[12] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM578 VSS WL0[12] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM579 VSS WL0[12] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM580 VSS WL0[12] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM581 VSS WL0[12] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM582 VSS WL0[12] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM583 VSS WL0[12] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM584 VSS WL0[12] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM585 VSS WL0[12] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM586 VSS WL0[12] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM587 VSS WL0[12] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM588 VSS WL0[12] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM589 VSS WL0[12] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM590 VSS WL0[12] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM591 VSS WL0[12] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM592 VSS WL0[12] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM593 VSS WL0[12] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM594 VSS WL0[12] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM595 VSS WL0[12] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM596 VSS WL0[12] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM597 VSS WL0[12] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM598 VSS WL0[12] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM599 VSS WL0[12] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM600 VSS WL0[12] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM601 VSS WL0[12] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM602 VSS WL0[12] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM603 VSS WL0[12] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM604 VSS WL0[12] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM605 VSS WL0[12] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM606 VSS WL0[12] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM607 VSS WL0[12] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM608 VSS WL0[12] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM609 VSS WL0[12] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM610 VSS WL0[12] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM611 VSS WL0[12] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM612 VSS WL0[12] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM613 VSS WL0[12] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM614 VSS WL0[12] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM615 VSS WL0[12] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM616 VSS WL0[12] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM617 VSS WL0[12] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM618 VSS WL0[12] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM619 VSS WL0[12] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM620 VSS WL0[12] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM621 VSS WL0[12] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM622 VSS WL0[12] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM623 VSS WL0[12] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM624 VSS WL0[12] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM625 VSS WL0[12] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM626 VSS WL0[12] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM627 VSS WL0[12] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM628 VSS WL0[12] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM629 VSS WL0[12] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM630 VSS WL0[12] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM631 VSS WL0[12] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0xd0
XM632 VSS WL0[13] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM633 VSS WL0[13] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM634 VSS WL0[13] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM635 VSS WL0[13] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM636 VSS WL0[13] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM637 VSS WL0[13] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM638 VSS WL0[13] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM639 VSS WL0[13] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM640 VSS WL0[13] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM641 VSS WL0[13] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM642 VSS WL0[13] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM643 VSS WL0[13] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM644 VSS WL0[13] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM645 VSS WL0[13] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM646 VSS WL0[13] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM647 VSS WL0[13] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM648 VSS WL0[13] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM649 VSS WL0[13] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM650 VSS WL0[13] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM651 VSS WL0[13] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM652 VSS WL0[13] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM653 VSS WL0[13] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM654 VSS WL0[13] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM655 VSS WL0[13] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM656 VSS WL0[13] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM657 VSS WL0[13] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM658 VSS WL0[13] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM659 VSS WL0[13] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM660 VSS WL0[13] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM661 VSS WL0[13] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM662 VSS WL0[13] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM663 VSS WL0[13] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM664 VSS WL0[13] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM665 VSS WL0[13] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM666 VSS WL0[13] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM667 VSS WL0[13] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM668 VSS WL0[13] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM669 VSS WL0[13] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM670 VSS WL0[13] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM671 VSS WL0[13] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM672 VSS WL0[13] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM673 VSS WL0[13] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM674 VSS WL0[13] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM675 VSS WL0[13] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM676 VSS WL0[13] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM677 VSS WL0[13] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM678 VSS WL0[13] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM679 VSS WL0[13] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM680 VSS WL0[13] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM681 VSS WL0[13] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM682 VSS WL0[13] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM683 VSS WL0[13] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0xe0
XM684 VSS WL0[14] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM685 VSS WL0[14] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM686 VSS WL0[14] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM687 VSS WL0[14] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM688 VSS WL0[14] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM689 VSS WL0[14] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM690 VSS WL0[14] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM691 VSS WL0[14] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM692 VSS WL0[14] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM693 VSS WL0[14] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM694 VSS WL0[14] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM695 VSS WL0[14] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM696 VSS WL0[14] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM697 VSS WL0[14] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM698 VSS WL0[14] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM699 VSS WL0[14] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM700 VSS WL0[14] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM701 VSS WL0[14] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM702 VSS WL0[14] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM703 VSS WL0[14] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM704 VSS WL0[14] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM705 VSS WL0[14] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM706 VSS WL0[14] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM707 VSS WL0[14] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM708 VSS WL0[14] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM709 VSS WL0[14] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM710 VSS WL0[14] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM711 VSS WL0[14] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM712 VSS WL0[14] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM713 VSS WL0[14] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM714 VSS WL0[14] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM715 VSS WL0[14] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM716 VSS WL0[14] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM717 VSS WL0[14] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM718 VSS WL0[14] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM719 VSS WL0[14] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM720 VSS WL0[14] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM721 VSS WL0[14] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM722 VSS WL0[14] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0xf0
XM723 VSS WL0[15] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM724 VSS WL0[15] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM725 VSS WL0[15] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM726 VSS WL0[15] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM727 VSS WL0[15] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM728 VSS WL0[15] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM729 VSS WL0[15] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM730 VSS WL0[15] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM731 VSS WL0[15] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM732 VSS WL0[15] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM733 VSS WL0[15] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM734 VSS WL0[15] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM735 VSS WL0[15] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM736 VSS WL0[15] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM737 VSS WL0[15] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM738 VSS WL0[15] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM739 VSS WL0[15] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM740 VSS WL0[15] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM741 VSS WL0[15] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM742 VSS WL0[15] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM743 VSS WL0[15] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM744 VSS WL0[15] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM745 VSS WL0[15] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM746 VSS WL0[15] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM747 VSS WL0[15] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM748 VSS WL0[15] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM749 VSS WL0[15] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM750 VSS WL0[15] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM751 VSS WL0[15] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM752 VSS WL0[15] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM753 VSS WL0[15] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM754 VSS WL0[15] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM755 VSS WL0[15] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM756 VSS WL0[15] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM757 VSS WL0[15] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM758 VSS WL0[15] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM759 VSS WL0[15] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM760 VSS WL0[15] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM761 VSS WL0[15] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM762 VSS WL0[15] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM763 VSS WL0[15] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM764 VSS WL0[15] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM765 VSS WL0[15] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM766 VSS WL0[15] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM767 VSS WL0[15] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM768 VSS WL0[15] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM769 VSS WL0[15] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM770 VSS WL0[15] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM771 VSS WL0[15] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM772 VSS WL0[15] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM773 VSS WL0[15] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x100
XM774 VSS WL0[16] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM775 VSS WL0[16] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM776 VSS WL0[16] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM777 VSS WL0[16] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM778 VSS WL0[16] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM779 VSS WL0[16] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM780 VSS WL0[16] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM781 VSS WL0[16] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM782 VSS WL0[16] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM783 VSS WL0[16] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM784 VSS WL0[16] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM785 VSS WL0[16] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM786 VSS WL0[16] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM787 VSS WL0[16] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM788 VSS WL0[16] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM789 VSS WL0[16] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM790 VSS WL0[16] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM791 VSS WL0[16] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM792 VSS WL0[16] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM793 VSS WL0[16] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM794 VSS WL0[16] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM795 VSS WL0[16] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM796 VSS WL0[16] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM797 VSS WL0[16] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM798 VSS WL0[16] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM799 VSS WL0[16] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM800 VSS WL0[16] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM801 VSS WL0[16] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM802 VSS WL0[16] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM803 VSS WL0[16] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM804 VSS WL0[16] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM805 VSS WL0[16] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM806 VSS WL0[16] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM807 VSS WL0[16] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM808 VSS WL0[16] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM809 VSS WL0[16] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM810 VSS WL0[16] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM811 VSS WL0[16] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM812 VSS WL0[16] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM813 VSS WL0[16] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM814 VSS WL0[16] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM815 VSS WL0[16] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM816 VSS WL0[16] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM817 VSS WL0[16] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM818 VSS WL0[16] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM819 VSS WL0[16] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM820 VSS WL0[16] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM821 VSS WL0[16] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM822 VSS WL0[16] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM823 VSS WL0[16] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM824 VSS WL0[16] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM825 VSS WL0[16] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM826 VSS WL0[16] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM827 VSS WL0[16] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM828 VSS WL0[16] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM829 VSS WL0[16] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM830 VSS WL0[16] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM831 VSS WL0[16] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM832 VSS WL0[16] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM833 VSS WL0[16] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x110
XM834 VSS WL0[17] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM835 VSS WL0[17] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM836 VSS WL0[17] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM837 VSS WL0[17] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM838 VSS WL0[17] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM839 VSS WL0[17] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM840 VSS WL0[17] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM841 VSS WL0[17] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM842 VSS WL0[17] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM843 VSS WL0[17] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM844 VSS WL0[17] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM845 VSS WL0[17] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM846 VSS WL0[17] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM847 VSS WL0[17] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM848 VSS WL0[17] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM849 VSS WL0[17] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM850 VSS WL0[17] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM851 VSS WL0[17] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM852 VSS WL0[17] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM853 VSS WL0[17] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM854 VSS WL0[17] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM855 VSS WL0[17] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM856 VSS WL0[17] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM857 VSS WL0[17] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM858 VSS WL0[17] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM859 VSS WL0[17] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM860 VSS WL0[17] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM861 VSS WL0[17] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM862 VSS WL0[17] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM863 VSS WL0[17] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM864 VSS WL0[17] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM865 VSS WL0[17] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM866 VSS WL0[17] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM867 VSS WL0[17] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM868 VSS WL0[17] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM869 VSS WL0[17] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM870 VSS WL0[17] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM871 VSS WL0[17] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM872 VSS WL0[17] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM873 VSS WL0[17] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM874 VSS WL0[17] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM875 VSS WL0[17] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x120
XM876 VSS WL0[18] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM877 VSS WL0[18] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM878 VSS WL0[18] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM879 VSS WL0[18] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM880 VSS WL0[18] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM881 VSS WL0[18] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM882 VSS WL0[18] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM883 VSS WL0[18] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM884 VSS WL0[18] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM885 VSS WL0[18] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM886 VSS WL0[18] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM887 VSS WL0[18] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM888 VSS WL0[18] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM889 VSS WL0[18] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM890 VSS WL0[18] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM891 VSS WL0[18] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM892 VSS WL0[18] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM893 VSS WL0[18] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM894 VSS WL0[18] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM895 VSS WL0[18] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM896 VSS WL0[18] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM897 VSS WL0[18] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM898 VSS WL0[18] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM899 VSS WL0[18] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM900 VSS WL0[18] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM901 VSS WL0[18] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM902 VSS WL0[18] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM903 VSS WL0[18] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM904 VSS WL0[18] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM905 VSS WL0[18] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM906 VSS WL0[18] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM907 VSS WL0[18] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM908 VSS WL0[18] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM909 VSS WL0[18] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM910 VSS WL0[18] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM911 VSS WL0[18] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM912 VSS WL0[18] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM913 VSS WL0[18] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM914 VSS WL0[18] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM915 VSS WL0[18] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM916 VSS WL0[18] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM917 VSS WL0[18] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM918 VSS WL0[18] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x130
XM919 VSS WL0[19] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM920 VSS WL0[19] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM921 VSS WL0[19] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM922 VSS WL0[19] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM923 VSS WL0[19] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM924 VSS WL0[19] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM925 VSS WL0[19] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM926 VSS WL0[19] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM927 VSS WL0[19] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM928 VSS WL0[19] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM929 VSS WL0[19] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM930 VSS WL0[19] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM931 VSS WL0[19] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM932 VSS WL0[19] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM933 VSS WL0[19] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM934 VSS WL0[19] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM935 VSS WL0[19] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM936 VSS WL0[19] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM937 VSS WL0[19] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM938 VSS WL0[19] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM939 VSS WL0[19] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM940 VSS WL0[19] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM941 VSS WL0[19] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM942 VSS WL0[19] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM943 VSS WL0[19] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM944 VSS WL0[19] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM945 VSS WL0[19] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM946 VSS WL0[19] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM947 VSS WL0[19] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM948 VSS WL0[19] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM949 VSS WL0[19] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM950 VSS WL0[19] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM951 VSS WL0[19] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM952 VSS WL0[19] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM953 VSS WL0[19] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM954 VSS WL0[19] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM955 VSS WL0[19] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM956 VSS WL0[19] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM957 VSS WL0[19] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM958 VSS WL0[19] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM959 VSS WL0[19] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM960 VSS WL0[19] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM961 VSS WL0[19] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM962 VSS WL0[19] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM963 VSS WL0[19] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM964 VSS WL0[19] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM965 VSS WL0[19] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM966 VSS WL0[19] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM967 VSS WL0[19] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM968 VSS WL0[19] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM969 VSS WL0[19] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM970 VSS WL0[19] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM971 VSS WL0[19] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM972 VSS WL0[19] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM973 VSS WL0[19] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM974 VSS WL0[19] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM975 VSS WL0[19] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM976 VSS WL0[19] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM977 VSS WL0[19] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM978 VSS WL0[19] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM979 VSS WL0[19] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM980 VSS WL0[19] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM981 VSS WL0[19] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x140
XM982 VSS WL0[20] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM983 VSS WL0[20] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM984 VSS WL0[20] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM985 VSS WL0[20] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM986 VSS WL0[20] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM987 VSS WL0[20] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM988 VSS WL0[20] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM989 VSS WL0[20] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM990 VSS WL0[20] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM991 VSS WL0[20] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM992 VSS WL0[20] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM993 VSS WL0[20] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM994 VSS WL0[20] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM995 VSS WL0[20] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM996 VSS WL0[20] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM997 VSS WL0[20] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM998 VSS WL0[20] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM999 VSS WL0[20] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1000 VSS WL0[20] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1001 VSS WL0[20] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1002 VSS WL0[20] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1003 VSS WL0[20] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1004 VSS WL0[20] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1005 VSS WL0[20] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1006 VSS WL0[20] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1007 VSS WL0[20] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1008 VSS WL0[20] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1009 VSS WL0[20] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1010 VSS WL0[20] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1011 VSS WL0[20] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1012 VSS WL0[20] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1013 VSS WL0[20] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1014 VSS WL0[20] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1015 VSS WL0[20] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1016 VSS WL0[20] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1017 VSS WL0[20] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1018 VSS WL0[20] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1019 VSS WL0[20] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1020 VSS WL0[20] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1021 VSS WL0[20] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1022 VSS WL0[20] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1023 VSS WL0[20] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1024 VSS WL0[20] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1025 VSS WL0[20] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1026 VSS WL0[20] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1027 VSS WL0[20] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1028 VSS WL0[20] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1029 VSS WL0[20] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1030 VSS WL0[20] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1031 VSS WL0[20] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1032 VSS WL0[20] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1033 VSS WL0[20] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1034 VSS WL0[20] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1035 VSS WL0[20] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1036 VSS WL0[20] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1037 VSS WL0[20] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x150
XM1038 VSS WL0[21] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1039 VSS WL0[21] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1040 VSS WL0[21] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1041 VSS WL0[21] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1042 VSS WL0[21] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1043 VSS WL0[21] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1044 VSS WL0[21] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1045 VSS WL0[21] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1046 VSS WL0[21] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1047 VSS WL0[21] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1048 VSS WL0[21] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1049 VSS WL0[21] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1050 VSS WL0[21] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1051 VSS WL0[21] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1052 VSS WL0[21] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1053 VSS WL0[21] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1054 VSS WL0[21] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1055 VSS WL0[21] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1056 VSS WL0[21] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1057 VSS WL0[21] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1058 VSS WL0[21] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1059 VSS WL0[21] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1060 VSS WL0[21] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1061 VSS WL0[21] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1062 VSS WL0[21] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1063 VSS WL0[21] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1064 VSS WL0[21] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1065 VSS WL0[21] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1066 VSS WL0[21] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1067 VSS WL0[21] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1068 VSS WL0[21] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1069 VSS WL0[21] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1070 VSS WL0[21] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1071 VSS WL0[21] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1072 VSS WL0[21] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1073 VSS WL0[21] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1074 VSS WL0[21] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1075 VSS WL0[21] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1076 VSS WL0[21] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1077 VSS WL0[21] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1078 VSS WL0[21] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1079 VSS WL0[21] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1080 VSS WL0[21] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1081 VSS WL0[21] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1082 VSS WL0[21] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1083 VSS WL0[21] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1084 VSS WL0[21] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1085 VSS WL0[21] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1086 VSS WL0[21] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1087 VSS WL0[21] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1088 VSS WL0[21] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1089 VSS WL0[21] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1090 VSS WL0[21] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1091 VSS WL0[21] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1092 VSS WL0[21] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1093 VSS WL0[21] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1094 VSS WL0[21] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1095 VSS WL0[21] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1096 VSS WL0[21] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1097 VSS WL0[21] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1098 VSS WL0[21] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1099 VSS WL0[21] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1100 VSS WL0[21] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1101 VSS WL0[21] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1102 VSS WL0[21] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1103 VSS WL0[21] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1104 VSS WL0[21] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1105 VSS WL0[21] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1106 VSS WL0[21] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1107 VSS WL0[21] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1108 VSS WL0[21] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1109 VSS WL0[21] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1110 VSS WL0[21] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1111 VSS WL0[21] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1112 VSS WL0[21] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1113 VSS WL0[21] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x160
XM1114 VSS WL0[22] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1115 VSS WL0[22] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1116 VSS WL0[22] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1117 VSS WL0[22] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1118 VSS WL0[22] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1119 VSS WL0[22] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1120 VSS WL0[22] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1121 VSS WL0[22] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1122 VSS WL0[22] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1123 VSS WL0[22] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1124 VSS WL0[22] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1125 VSS WL0[22] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1126 VSS WL0[22] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1127 VSS WL0[22] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1128 VSS WL0[22] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1129 VSS WL0[22] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1130 VSS WL0[22] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1131 VSS WL0[22] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1132 VSS WL0[22] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1133 VSS WL0[22] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1134 VSS WL0[22] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1135 VSS WL0[22] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1136 VSS WL0[22] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1137 VSS WL0[22] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1138 VSS WL0[22] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1139 VSS WL0[22] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1140 VSS WL0[22] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1141 VSS WL0[22] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1142 VSS WL0[22] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1143 VSS WL0[22] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1144 VSS WL0[22] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1145 VSS WL0[22] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1146 VSS WL0[22] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1147 VSS WL0[22] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1148 VSS WL0[22] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1149 VSS WL0[22] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1150 VSS WL0[22] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1151 VSS WL0[22] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1152 VSS WL0[22] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1153 VSS WL0[22] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1154 VSS WL0[22] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1155 VSS WL0[22] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1156 VSS WL0[22] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1157 VSS WL0[22] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1158 VSS WL0[22] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1159 VSS WL0[22] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1160 VSS WL0[22] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1161 VSS WL0[22] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1162 VSS WL0[22] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1163 VSS WL0[22] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1164 VSS WL0[22] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1165 VSS WL0[22] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1166 VSS WL0[22] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x170
XM1167 VSS WL0[23] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1168 VSS WL0[23] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1169 VSS WL0[23] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1170 VSS WL0[23] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1171 VSS WL0[23] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1172 VSS WL0[23] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1173 VSS WL0[23] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1174 VSS WL0[23] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1175 VSS WL0[23] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1176 VSS WL0[23] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1177 VSS WL0[23] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1178 VSS WL0[23] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1179 VSS WL0[23] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1180 VSS WL0[23] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1181 VSS WL0[23] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1182 VSS WL0[23] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1183 VSS WL0[23] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1184 VSS WL0[23] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1185 VSS WL0[23] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1186 VSS WL0[23] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1187 VSS WL0[23] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1188 VSS WL0[23] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1189 VSS WL0[23] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1190 VSS WL0[23] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1191 VSS WL0[23] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1192 VSS WL0[23] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1193 VSS WL0[23] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1194 VSS WL0[23] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1195 VSS WL0[23] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1196 VSS WL0[23] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1197 VSS WL0[23] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1198 VSS WL0[23] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1199 VSS WL0[23] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1200 VSS WL0[23] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1201 VSS WL0[23] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1202 VSS WL0[23] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1203 VSS WL0[23] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1204 VSS WL0[23] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1205 VSS WL0[23] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1206 VSS WL0[23] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1207 VSS WL0[23] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1208 VSS WL0[23] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1209 VSS WL0[23] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1210 VSS WL0[23] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1211 VSS WL0[23] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1212 VSS WL0[23] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1213 VSS WL0[23] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1214 VSS WL0[23] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1215 VSS WL0[23] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1216 VSS WL0[23] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1217 VSS WL0[23] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1218 VSS WL0[23] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1219 VSS WL0[23] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1220 VSS WL0[23] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1221 VSS WL0[23] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1222 VSS WL0[23] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1223 VSS WL0[23] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1224 VSS WL0[23] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1225 VSS WL0[23] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x180
XM1226 VSS WL0[24] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1227 VSS WL0[24] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1228 VSS WL0[24] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1229 VSS WL0[24] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1230 VSS WL0[24] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1231 VSS WL0[24] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1232 VSS WL0[24] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1233 VSS WL0[24] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1234 VSS WL0[24] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1235 VSS WL0[24] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1236 VSS WL0[24] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1237 VSS WL0[24] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1238 VSS WL0[24] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1239 VSS WL0[24] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1240 VSS WL0[24] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1241 VSS WL0[24] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1242 VSS WL0[24] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1243 VSS WL0[24] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1244 VSS WL0[24] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1245 VSS WL0[24] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1246 VSS WL0[24] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1247 VSS WL0[24] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1248 VSS WL0[24] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1249 VSS WL0[24] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1250 VSS WL0[24] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1251 VSS WL0[24] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1252 VSS WL0[24] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1253 VSS WL0[24] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1254 VSS WL0[24] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1255 VSS WL0[24] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1256 VSS WL0[24] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1257 VSS WL0[24] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1258 VSS WL0[24] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1259 VSS WL0[24] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1260 VSS WL0[24] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1261 VSS WL0[24] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1262 VSS WL0[24] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1263 VSS WL0[24] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1264 VSS WL0[24] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1265 VSS WL0[24] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1266 VSS WL0[24] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1267 VSS WL0[24] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1268 VSS WL0[24] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1269 VSS WL0[24] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1270 VSS WL0[24] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1271 VSS WL0[24] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1272 VSS WL0[24] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1273 VSS WL0[24] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1274 VSS WL0[24] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1275 VSS WL0[24] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1276 VSS WL0[24] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1277 VSS WL0[24] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1278 VSS WL0[24] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1279 VSS WL0[24] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1280 VSS WL0[24] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1281 VSS WL0[24] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1282 VSS WL0[24] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1283 VSS WL0[24] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1284 VSS WL0[24] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1285 VSS WL0[24] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1286 VSS WL0[24] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1287 VSS WL0[24] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1288 VSS WL0[24] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1289 VSS WL0[24] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1290 VSS WL0[24] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1291 VSS WL0[24] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1292 VSS WL0[24] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1293 VSS WL0[24] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1294 VSS WL0[24] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1295 VSS WL0[24] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1296 VSS WL0[24] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1297 VSS WL0[24] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1298 VSS WL0[24] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1299 VSS WL0[24] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1300 VSS WL0[24] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x190
XM1301 VSS WL0[25] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1302 VSS WL0[25] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1303 VSS WL0[25] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1304 VSS WL0[25] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1305 VSS WL0[25] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1306 VSS WL0[25] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1307 VSS WL0[25] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1308 VSS WL0[25] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1309 VSS WL0[25] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1310 VSS WL0[25] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1311 VSS WL0[25] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1312 VSS WL0[25] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1313 VSS WL0[25] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1314 VSS WL0[25] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1315 VSS WL0[25] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1316 VSS WL0[25] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1317 VSS WL0[25] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1318 VSS WL0[25] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1319 VSS WL0[25] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1320 VSS WL0[25] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1321 VSS WL0[25] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1322 VSS WL0[25] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1323 VSS WL0[25] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1324 VSS WL0[25] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1325 VSS WL0[25] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1326 VSS WL0[25] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1327 VSS WL0[25] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1328 VSS WL0[25] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1329 VSS WL0[25] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1330 VSS WL0[25] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1331 VSS WL0[25] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1332 VSS WL0[25] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1333 VSS WL0[25] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1334 VSS WL0[25] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1335 VSS WL0[25] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1336 VSS WL0[25] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1337 VSS WL0[25] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1338 VSS WL0[25] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1339 VSS WL0[25] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1340 VSS WL0[25] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1341 VSS WL0[25] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1342 VSS WL0[25] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1343 VSS WL0[25] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1344 VSS WL0[25] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1345 VSS WL0[25] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1346 VSS WL0[25] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x1a0
XM1347 VSS WL0[26] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1348 VSS WL0[26] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1349 VSS WL0[26] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1350 VSS WL0[26] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1351 VSS WL0[26] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1352 VSS WL0[26] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1353 VSS WL0[26] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1354 VSS WL0[26] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1355 VSS WL0[26] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1356 VSS WL0[26] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1357 VSS WL0[26] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1358 VSS WL0[26] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1359 VSS WL0[26] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1360 VSS WL0[26] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1361 VSS WL0[26] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1362 VSS WL0[26] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1363 VSS WL0[26] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1364 VSS WL0[26] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1365 VSS WL0[26] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1366 VSS WL0[26] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1367 VSS WL0[26] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1368 VSS WL0[26] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1369 VSS WL0[26] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1370 VSS WL0[26] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1371 VSS WL0[26] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1372 VSS WL0[26] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1373 VSS WL0[26] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1374 VSS WL0[26] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1375 VSS WL0[26] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1376 VSS WL0[26] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1377 VSS WL0[26] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1378 VSS WL0[26] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1379 VSS WL0[26] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1380 VSS WL0[26] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1381 VSS WL0[26] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1382 VSS WL0[26] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1383 VSS WL0[26] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1384 VSS WL0[26] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1385 VSS WL0[26] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1386 VSS WL0[26] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1387 VSS WL0[26] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1388 VSS WL0[26] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1389 VSS WL0[26] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1390 VSS WL0[26] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1391 VSS WL0[26] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1392 VSS WL0[26] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1393 VSS WL0[26] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1394 VSS WL0[26] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1395 VSS WL0[26] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1396 VSS WL0[26] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1397 VSS WL0[26] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1398 VSS WL0[26] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1399 VSS WL0[26] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1400 VSS WL0[26] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x1b0
XM1401 VSS WL0[27] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1402 VSS WL0[27] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1403 VSS WL0[27] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1404 VSS WL0[27] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1405 VSS WL0[27] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1406 VSS WL0[27] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1407 VSS WL0[27] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1408 VSS WL0[27] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1409 VSS WL0[27] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1410 VSS WL0[27] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1411 VSS WL0[27] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1412 VSS WL0[27] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1413 VSS WL0[27] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1414 VSS WL0[27] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1415 VSS WL0[27] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1416 VSS WL0[27] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1417 VSS WL0[27] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1418 VSS WL0[27] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1419 VSS WL0[27] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1420 VSS WL0[27] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1421 VSS WL0[27] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1422 VSS WL0[27] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1423 VSS WL0[27] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1424 VSS WL0[27] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1425 VSS WL0[27] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1426 VSS WL0[27] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1427 VSS WL0[27] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1428 VSS WL0[27] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1429 VSS WL0[27] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1430 VSS WL0[27] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1431 VSS WL0[27] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1432 VSS WL0[27] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1433 VSS WL0[27] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1434 VSS WL0[27] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1435 VSS WL0[27] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1436 VSS WL0[27] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1437 VSS WL0[27] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1438 VSS WL0[27] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1439 VSS WL0[27] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1440 VSS WL0[27] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1441 VSS WL0[27] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1442 VSS WL0[27] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1443 VSS WL0[27] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1444 VSS WL0[27] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1445 VSS WL0[27] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1446 VSS WL0[27] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1447 VSS WL0[27] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1448 VSS WL0[27] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1449 VSS WL0[27] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1450 VSS WL0[27] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1451 VSS WL0[27] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1452 VSS WL0[27] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x1c0
XM1453 VSS WL0[28] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1454 VSS WL0[28] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1455 VSS WL0[28] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1456 VSS WL0[28] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1457 VSS WL0[28] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1458 VSS WL0[28] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1459 VSS WL0[28] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1460 VSS WL0[28] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1461 VSS WL0[28] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1462 VSS WL0[28] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1463 VSS WL0[28] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1464 VSS WL0[28] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1465 VSS WL0[28] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1466 VSS WL0[28] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1467 VSS WL0[28] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1468 VSS WL0[28] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1469 VSS WL0[28] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1470 VSS WL0[28] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1471 VSS WL0[28] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1472 VSS WL0[28] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1473 VSS WL0[28] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1474 VSS WL0[28] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1475 VSS WL0[28] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1476 VSS WL0[28] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1477 VSS WL0[28] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1478 VSS WL0[28] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1479 VSS WL0[28] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1480 VSS WL0[28] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1481 VSS WL0[28] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1482 VSS WL0[28] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1483 VSS WL0[28] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1484 VSS WL0[28] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1485 VSS WL0[28] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1486 VSS WL0[28] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1487 VSS WL0[28] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x1d0
XM1488 VSS WL0[29] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1489 VSS WL0[29] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1490 VSS WL0[29] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1491 VSS WL0[29] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1492 VSS WL0[29] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1493 VSS WL0[29] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1494 VSS WL0[29] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1495 VSS WL0[29] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1496 VSS WL0[29] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1497 VSS WL0[29] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1498 VSS WL0[29] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1499 VSS WL0[29] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1500 VSS WL0[29] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1501 VSS WL0[29] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1502 VSS WL0[29] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1503 VSS WL0[29] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1504 VSS WL0[29] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1505 VSS WL0[29] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1506 VSS WL0[29] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1507 VSS WL0[29] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1508 VSS WL0[29] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1509 VSS WL0[29] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1510 VSS WL0[29] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1511 VSS WL0[29] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1512 VSS WL0[29] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1513 VSS WL0[29] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1514 VSS WL0[29] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1515 VSS WL0[29] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1516 VSS WL0[29] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1517 VSS WL0[29] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1518 VSS WL0[29] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1519 VSS WL0[29] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1520 VSS WL0[29] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1521 VSS WL0[29] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1522 VSS WL0[29] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1523 VSS WL0[29] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1524 VSS WL0[29] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1525 VSS WL0[29] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1526 VSS WL0[29] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1527 VSS WL0[29] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1528 VSS WL0[29] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1529 VSS WL0[29] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1530 VSS WL0[29] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1531 VSS WL0[29] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1532 VSS WL0[29] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1533 VSS WL0[29] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1534 VSS WL0[29] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1535 VSS WL0[29] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1536 VSS WL0[29] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1537 VSS WL0[29] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1538 VSS WL0[29] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1539 VSS WL0[29] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x1e0
XM1540 VSS WL0[30] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1541 VSS WL0[30] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1542 VSS WL0[30] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1543 VSS WL0[30] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1544 VSS WL0[30] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1545 VSS WL0[30] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1546 VSS WL0[30] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1547 VSS WL0[30] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1548 VSS WL0[30] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1549 VSS WL0[30] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1550 VSS WL0[30] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1551 VSS WL0[30] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1552 VSS WL0[30] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1553 VSS WL0[30] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1554 VSS WL0[30] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1555 VSS WL0[30] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1556 VSS WL0[30] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1557 VSS WL0[30] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1558 VSS WL0[30] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1559 VSS WL0[30] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1560 VSS WL0[30] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1561 VSS WL0[30] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1562 VSS WL0[30] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1563 VSS WL0[30] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1564 VSS WL0[30] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1565 VSS WL0[30] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1566 VSS WL0[30] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1567 VSS WL0[30] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1568 VSS WL0[30] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1569 VSS WL0[30] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1570 VSS WL0[30] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1571 VSS WL0[30] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1572 VSS WL0[30] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1573 VSS WL0[30] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1574 VSS WL0[30] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1575 VSS WL0[30] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1576 VSS WL0[30] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1577 VSS WL0[30] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1578 VSS WL0[30] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1579 VSS WL0[30] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1580 VSS WL0[30] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1581 VSS WL0[30] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1582 VSS WL0[30] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1583 VSS WL0[30] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1584 VSS WL0[30] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x1f0
XM1585 VSS WL0[31] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1586 VSS WL0[31] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1587 VSS WL0[31] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1588 VSS WL0[31] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1589 VSS WL0[31] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1590 VSS WL0[31] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1591 VSS WL0[31] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1592 VSS WL0[31] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1593 VSS WL0[31] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1594 VSS WL0[31] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1595 VSS WL0[31] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1596 VSS WL0[31] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1597 VSS WL0[31] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1598 VSS WL0[31] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1599 VSS WL0[31] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1600 VSS WL0[31] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1601 VSS WL0[31] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1602 VSS WL0[31] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1603 VSS WL0[31] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1604 VSS WL0[31] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1605 VSS WL0[31] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1606 VSS WL0[31] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1607 VSS WL0[31] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1608 VSS WL0[31] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1609 VSS WL0[31] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1610 VSS WL0[31] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1611 VSS WL0[31] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1612 VSS WL0[31] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1613 VSS WL0[31] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1614 VSS WL0[31] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1615 VSS WL0[31] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1616 VSS WL0[31] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1617 VSS WL0[31] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1618 VSS WL0[31] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1619 VSS WL0[31] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1620 VSS WL0[31] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1621 VSS WL0[31] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1622 VSS WL0[31] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1623 VSS WL0[31] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1624 VSS WL0[31] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1625 VSS WL0[31] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1626 VSS WL0[31] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1627 VSS WL0[31] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1628 VSS WL0[31] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1629 VSS WL0[31] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1630 VSS WL0[31] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1631 VSS WL0[31] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1632 VSS WL0[31] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x200
XM1633 VSS WL0[32] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1634 VSS WL0[32] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1635 VSS WL0[32] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1636 VSS WL0[32] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1637 VSS WL0[32] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1638 VSS WL0[32] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1639 VSS WL0[32] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1640 VSS WL0[32] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1641 VSS WL0[32] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1642 VSS WL0[32] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1643 VSS WL0[32] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1644 VSS WL0[32] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1645 VSS WL0[32] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1646 VSS WL0[32] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1647 VSS WL0[32] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1648 VSS WL0[32] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1649 VSS WL0[32] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1650 VSS WL0[32] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1651 VSS WL0[32] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1652 VSS WL0[32] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1653 VSS WL0[32] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1654 VSS WL0[32] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1655 VSS WL0[32] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1656 VSS WL0[32] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1657 VSS WL0[32] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1658 VSS WL0[32] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1659 VSS WL0[32] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1660 VSS WL0[32] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1661 VSS WL0[32] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1662 VSS WL0[32] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1663 VSS WL0[32] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1664 VSS WL0[32] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1665 VSS WL0[32] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1666 VSS WL0[32] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1667 VSS WL0[32] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1668 VSS WL0[32] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1669 VSS WL0[32] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1670 VSS WL0[32] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1671 VSS WL0[32] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1672 VSS WL0[32] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1673 VSS WL0[32] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1674 VSS WL0[32] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1675 VSS WL0[32] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1676 VSS WL0[32] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1677 VSS WL0[32] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1678 VSS WL0[32] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1679 VSS WL0[32] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1680 VSS WL0[32] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1681 VSS WL0[32] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1682 VSS WL0[32] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x210
XM1683 VSS WL0[33] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1684 VSS WL0[33] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1685 VSS WL0[33] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1686 VSS WL0[33] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1687 VSS WL0[33] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1688 VSS WL0[33] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1689 VSS WL0[33] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1690 VSS WL0[33] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1691 VSS WL0[33] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1692 VSS WL0[33] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1693 VSS WL0[33] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1694 VSS WL0[33] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1695 VSS WL0[33] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1696 VSS WL0[33] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1697 VSS WL0[33] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1698 VSS WL0[33] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1699 VSS WL0[33] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1700 VSS WL0[33] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1701 VSS WL0[33] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1702 VSS WL0[33] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1703 VSS WL0[33] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1704 VSS WL0[33] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1705 VSS WL0[33] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1706 VSS WL0[33] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1707 VSS WL0[33] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1708 VSS WL0[33] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1709 VSS WL0[33] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1710 VSS WL0[33] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1711 VSS WL0[33] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1712 VSS WL0[33] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1713 VSS WL0[33] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1714 VSS WL0[33] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1715 VSS WL0[33] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1716 VSS WL0[33] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1717 VSS WL0[33] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1718 VSS WL0[33] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1719 VSS WL0[33] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1720 VSS WL0[33] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1721 VSS WL0[33] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1722 VSS WL0[33] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1723 VSS WL0[33] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x220
XM1724 VSS WL0[34] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1725 VSS WL0[34] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1726 VSS WL0[34] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1727 VSS WL0[34] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1728 VSS WL0[34] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1729 VSS WL0[34] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1730 VSS WL0[34] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1731 VSS WL0[34] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1732 VSS WL0[34] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1733 VSS WL0[34] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1734 VSS WL0[34] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1735 VSS WL0[34] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1736 VSS WL0[34] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1737 VSS WL0[34] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1738 VSS WL0[34] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1739 VSS WL0[34] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1740 VSS WL0[34] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1741 VSS WL0[34] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1742 VSS WL0[34] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1743 VSS WL0[34] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1744 VSS WL0[34] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1745 VSS WL0[34] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1746 VSS WL0[34] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1747 VSS WL0[34] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1748 VSS WL0[34] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1749 VSS WL0[34] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1750 VSS WL0[34] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1751 VSS WL0[34] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1752 VSS WL0[34] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1753 VSS WL0[34] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1754 VSS WL0[34] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1755 VSS WL0[34] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1756 VSS WL0[34] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1757 VSS WL0[34] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1758 VSS WL0[34] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1759 VSS WL0[34] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1760 VSS WL0[34] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1761 VSS WL0[34] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1762 VSS WL0[34] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1763 VSS WL0[34] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1764 VSS WL0[34] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x230
XM1765 VSS WL0[35] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1766 VSS WL0[35] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1767 VSS WL0[35] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1768 VSS WL0[35] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1769 VSS WL0[35] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1770 VSS WL0[35] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1771 VSS WL0[35] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1772 VSS WL0[35] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1773 VSS WL0[35] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1774 VSS WL0[35] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1775 VSS WL0[35] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1776 VSS WL0[35] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1777 VSS WL0[35] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1778 VSS WL0[35] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1779 VSS WL0[35] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1780 VSS WL0[35] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1781 VSS WL0[35] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1782 VSS WL0[35] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1783 VSS WL0[35] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1784 VSS WL0[35] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1785 VSS WL0[35] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1786 VSS WL0[35] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1787 VSS WL0[35] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1788 VSS WL0[35] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1789 VSS WL0[35] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1790 VSS WL0[35] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1791 VSS WL0[35] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1792 VSS WL0[35] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1793 VSS WL0[35] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1794 VSS WL0[35] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1795 VSS WL0[35] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1796 VSS WL0[35] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1797 VSS WL0[35] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1798 VSS WL0[35] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1799 VSS WL0[35] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1800 VSS WL0[35] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1801 VSS WL0[35] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1802 VSS WL0[35] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1803 VSS WL0[35] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1804 VSS WL0[35] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1805 VSS WL0[35] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1806 VSS WL0[35] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1807 VSS WL0[35] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1808 VSS WL0[35] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x240
XM1809 VSS WL0[36] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1810 VSS WL0[36] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1811 VSS WL0[36] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1812 VSS WL0[36] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1813 VSS WL0[36] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1814 VSS WL0[36] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1815 VSS WL0[36] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1816 VSS WL0[36] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1817 VSS WL0[36] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1818 VSS WL0[36] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1819 VSS WL0[36] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1820 VSS WL0[36] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1821 VSS WL0[36] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1822 VSS WL0[36] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1823 VSS WL0[36] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1824 VSS WL0[36] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1825 VSS WL0[36] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1826 VSS WL0[36] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1827 VSS WL0[36] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1828 VSS WL0[36] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1829 VSS WL0[36] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1830 VSS WL0[36] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1831 VSS WL0[36] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1832 VSS WL0[36] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1833 VSS WL0[36] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1834 VSS WL0[36] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1835 VSS WL0[36] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1836 VSS WL0[36] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1837 VSS WL0[36] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1838 VSS WL0[36] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1839 VSS WL0[36] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1840 VSS WL0[36] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1841 VSS WL0[36] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1842 VSS WL0[36] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1843 VSS WL0[36] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1844 VSS WL0[36] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1845 VSS WL0[36] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1846 VSS WL0[36] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1847 VSS WL0[36] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1848 VSS WL0[36] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1849 VSS WL0[36] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1850 VSS WL0[36] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1851 VSS WL0[36] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1852 VSS WL0[36] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x250
XM1853 VSS WL0[37] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1854 VSS WL0[37] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1855 VSS WL0[37] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1856 VSS WL0[37] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1857 VSS WL0[37] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1858 VSS WL0[37] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1859 VSS WL0[37] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1860 VSS WL0[37] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1861 VSS WL0[37] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1862 VSS WL0[37] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1863 VSS WL0[37] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1864 VSS WL0[37] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1865 VSS WL0[37] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1866 VSS WL0[37] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1867 VSS WL0[37] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1868 VSS WL0[37] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1869 VSS WL0[37] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1870 VSS WL0[37] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1871 VSS WL0[37] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1872 VSS WL0[37] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1873 VSS WL0[37] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1874 VSS WL0[37] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1875 VSS WL0[37] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1876 VSS WL0[37] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1877 VSS WL0[37] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1878 VSS WL0[37] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1879 VSS WL0[37] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1880 VSS WL0[37] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1881 VSS WL0[37] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1882 VSS WL0[37] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1883 VSS WL0[37] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1884 VSS WL0[37] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1885 VSS WL0[37] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1886 VSS WL0[37] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1887 VSS WL0[37] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1888 VSS WL0[37] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1889 VSS WL0[37] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1890 VSS WL0[37] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1891 VSS WL0[37] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1892 VSS WL0[37] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1893 VSS WL0[37] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1894 VSS WL0[37] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1895 VSS WL0[37] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1896 VSS WL0[37] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1897 VSS WL0[37] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1898 VSS WL0[37] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1899 VSS WL0[37] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1900 VSS WL0[37] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1901 VSS WL0[37] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1902 VSS WL0[37] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1903 VSS WL0[37] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x260
XM1904 VSS WL0[38] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1905 VSS WL0[38] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1906 VSS WL0[38] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1907 VSS WL0[38] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1908 VSS WL0[38] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1909 VSS WL0[38] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1910 VSS WL0[38] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1911 VSS WL0[38] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1912 VSS WL0[38] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1913 VSS WL0[38] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1914 VSS WL0[38] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1915 VSS WL0[38] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1916 VSS WL0[38] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1917 VSS WL0[38] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1918 VSS WL0[38] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1919 VSS WL0[38] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1920 VSS WL0[38] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1921 VSS WL0[38] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1922 VSS WL0[38] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1923 VSS WL0[38] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1924 VSS WL0[38] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1925 VSS WL0[38] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1926 VSS WL0[38] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1927 VSS WL0[38] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1928 VSS WL0[38] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1929 VSS WL0[38] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1930 VSS WL0[38] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1931 VSS WL0[38] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1932 VSS WL0[38] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1933 VSS WL0[38] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1934 VSS WL0[38] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1935 VSS WL0[38] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1936 VSS WL0[38] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1937 VSS WL0[38] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1938 VSS WL0[38] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1939 VSS WL0[38] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x270
XM1940 VSS WL0[39] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1941 VSS WL0[39] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1942 VSS WL0[39] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1943 VSS WL0[39] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1944 VSS WL0[39] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1945 VSS WL0[39] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1946 VSS WL0[39] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1947 VSS WL0[39] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1948 VSS WL0[39] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1949 VSS WL0[39] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1950 VSS WL0[39] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1951 VSS WL0[39] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1952 VSS WL0[39] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1953 VSS WL0[39] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1954 VSS WL0[39] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1955 VSS WL0[39] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1956 VSS WL0[39] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1957 VSS WL0[39] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1958 VSS WL0[39] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1959 VSS WL0[39] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1960 VSS WL0[39] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1961 VSS WL0[39] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1962 VSS WL0[39] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1963 VSS WL0[39] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1964 VSS WL0[39] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1965 VSS WL0[39] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1966 VSS WL0[39] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1967 VSS WL0[39] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1968 VSS WL0[39] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1969 VSS WL0[39] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1970 VSS WL0[39] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1971 VSS WL0[39] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1972 VSS WL0[39] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1973 VSS WL0[39] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1974 VSS WL0[39] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1975 VSS WL0[39] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1976 VSS WL0[39] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1977 VSS WL0[39] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1978 VSS WL0[39] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1979 VSS WL0[39] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1980 VSS WL0[39] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1981 VSS WL0[39] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1982 VSS WL0[39] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1983 VSS WL0[39] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1984 VSS WL0[39] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1985 VSS WL0[39] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1986 VSS WL0[39] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1987 VSS WL0[39] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1988 VSS WL0[39] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1989 VSS WL0[39] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1990 VSS WL0[39] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1991 VSS WL0[39] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1992 VSS WL0[39] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1993 VSS WL0[39] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1994 VSS WL0[39] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1995 VSS WL0[39] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1996 VSS WL0[39] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1997 VSS WL0[39] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1998 VSS WL0[39] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM1999 VSS WL0[39] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2000 VSS WL0[39] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2001 VSS WL0[39] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2002 VSS WL0[39] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2003 VSS WL0[39] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2004 VSS WL0[39] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2005 VSS WL0[39] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2006 VSS WL0[39] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2007 VSS WL0[39] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x280
XM2008 VSS WL0[40] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2009 VSS WL0[40] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2010 VSS WL0[40] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2011 VSS WL0[40] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2012 VSS WL0[40] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2013 VSS WL0[40] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2014 VSS WL0[40] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2015 VSS WL0[40] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2016 VSS WL0[40] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2017 VSS WL0[40] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2018 VSS WL0[40] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2019 VSS WL0[40] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2020 VSS WL0[40] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2021 VSS WL0[40] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2022 VSS WL0[40] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2023 VSS WL0[40] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2024 VSS WL0[40] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2025 VSS WL0[40] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2026 VSS WL0[40] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2027 VSS WL0[40] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2028 VSS WL0[40] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2029 VSS WL0[40] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2030 VSS WL0[40] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2031 VSS WL0[40] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2032 VSS WL0[40] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2033 VSS WL0[40] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2034 VSS WL0[40] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2035 VSS WL0[40] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2036 VSS WL0[40] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2037 VSS WL0[40] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2038 VSS WL0[40] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2039 VSS WL0[40] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2040 VSS WL0[40] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2041 VSS WL0[40] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2042 VSS WL0[40] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2043 VSS WL0[40] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2044 VSS WL0[40] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2045 VSS WL0[40] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2046 VSS WL0[40] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2047 VSS WL0[40] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2048 VSS WL0[40] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2049 VSS WL0[40] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2050 VSS WL0[40] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2051 VSS WL0[40] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2052 VSS WL0[40] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2053 VSS WL0[40] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2054 VSS WL0[40] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2055 VSS WL0[40] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2056 VSS WL0[40] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2057 VSS WL0[40] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2058 VSS WL0[40] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x290
XM2059 VSS WL0[41] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2060 VSS WL0[41] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2061 VSS WL0[41] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2062 VSS WL0[41] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2063 VSS WL0[41] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2064 VSS WL0[41] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2065 VSS WL0[41] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2066 VSS WL0[41] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2067 VSS WL0[41] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2068 VSS WL0[41] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2069 VSS WL0[41] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2070 VSS WL0[41] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2071 VSS WL0[41] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2072 VSS WL0[41] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2073 VSS WL0[41] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2074 VSS WL0[41] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2075 VSS WL0[41] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2076 VSS WL0[41] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2077 VSS WL0[41] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2078 VSS WL0[41] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2079 VSS WL0[41] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2080 VSS WL0[41] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2081 VSS WL0[41] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2082 VSS WL0[41] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2083 VSS WL0[41] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2084 VSS WL0[41] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2085 VSS WL0[41] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2086 VSS WL0[41] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2087 VSS WL0[41] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2088 VSS WL0[41] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2089 VSS WL0[41] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2090 VSS WL0[41] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2091 VSS WL0[41] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2092 VSS WL0[41] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2093 VSS WL0[41] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2094 VSS WL0[41] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2095 VSS WL0[41] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2096 VSS WL0[41] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2097 VSS WL0[41] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2098 VSS WL0[41] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2099 VSS WL0[41] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2100 VSS WL0[41] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2101 VSS WL0[41] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2102 VSS WL0[41] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2103 VSS WL0[41] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2104 VSS WL0[41] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x2a0
XM2105 VSS WL0[42] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2106 VSS WL0[42] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2107 VSS WL0[42] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2108 VSS WL0[42] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2109 VSS WL0[42] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2110 VSS WL0[42] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2111 VSS WL0[42] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2112 VSS WL0[42] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2113 VSS WL0[42] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2114 VSS WL0[42] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2115 VSS WL0[42] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2116 VSS WL0[42] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2117 VSS WL0[42] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2118 VSS WL0[42] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2119 VSS WL0[42] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2120 VSS WL0[42] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2121 VSS WL0[42] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2122 VSS WL0[42] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2123 VSS WL0[42] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2124 VSS WL0[42] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2125 VSS WL0[42] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2126 VSS WL0[42] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2127 VSS WL0[42] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2128 VSS WL0[42] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2129 VSS WL0[42] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2130 VSS WL0[42] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2131 VSS WL0[42] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2132 VSS WL0[42] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2133 VSS WL0[42] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2134 VSS WL0[42] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2135 VSS WL0[42] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2136 VSS WL0[42] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2137 VSS WL0[42] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2138 VSS WL0[42] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2139 VSS WL0[42] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2140 VSS WL0[42] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2141 VSS WL0[42] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2142 VSS WL0[42] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2143 VSS WL0[42] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2144 VSS WL0[42] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2145 VSS WL0[42] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2146 VSS WL0[42] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2147 VSS WL0[42] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2148 VSS WL0[42] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2149 VSS WL0[42] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2150 VSS WL0[42] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2151 VSS WL0[42] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2152 VSS WL0[42] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2153 VSS WL0[42] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2154 VSS WL0[42] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2155 VSS WL0[42] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2156 VSS WL0[42] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2157 VSS WL0[42] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2158 VSS WL0[42] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2159 VSS WL0[42] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2160 VSS WL0[42] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2161 VSS WL0[42] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2162 VSS WL0[42] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2163 VSS WL0[42] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2164 VSS WL0[42] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x2b0
XM2165 VSS WL0[43] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2166 VSS WL0[43] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2167 VSS WL0[43] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2168 VSS WL0[43] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2169 VSS WL0[43] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2170 VSS WL0[43] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2171 VSS WL0[43] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2172 VSS WL0[43] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2173 VSS WL0[43] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2174 VSS WL0[43] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2175 VSS WL0[43] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2176 VSS WL0[43] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2177 VSS WL0[43] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2178 VSS WL0[43] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2179 VSS WL0[43] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2180 VSS WL0[43] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2181 VSS WL0[43] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2182 VSS WL0[43] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2183 VSS WL0[43] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2184 VSS WL0[43] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2185 VSS WL0[43] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2186 VSS WL0[43] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2187 VSS WL0[43] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2188 VSS WL0[43] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2189 VSS WL0[43] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2190 VSS WL0[43] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2191 VSS WL0[43] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2192 VSS WL0[43] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2193 VSS WL0[43] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2194 VSS WL0[43] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2195 VSS WL0[43] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2196 VSS WL0[43] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2197 VSS WL0[43] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2198 VSS WL0[43] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2199 VSS WL0[43] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2200 VSS WL0[43] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2201 VSS WL0[43] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2202 VSS WL0[43] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2203 VSS WL0[43] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2204 VSS WL0[43] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2205 VSS WL0[43] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2206 VSS WL0[43] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2207 VSS WL0[43] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2208 VSS WL0[43] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2209 VSS WL0[43] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2210 VSS WL0[43] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2211 VSS WL0[43] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2212 VSS WL0[43] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2213 VSS WL0[43] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2214 VSS WL0[43] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2215 VSS WL0[43] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2216 VSS WL0[43] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2217 VSS WL0[43] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2218 VSS WL0[43] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2219 VSS WL0[43] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2220 VSS WL0[43] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2221 VSS WL0[43] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2222 VSS WL0[43] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x2c0
XM2223 VSS WL0[44] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2224 VSS WL0[44] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2225 VSS WL0[44] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2226 VSS WL0[44] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2227 VSS WL0[44] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2228 VSS WL0[44] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2229 VSS WL0[44] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2230 VSS WL0[44] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2231 VSS WL0[44] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2232 VSS WL0[44] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2233 VSS WL0[44] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2234 VSS WL0[44] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2235 VSS WL0[44] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2236 VSS WL0[44] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2237 VSS WL0[44] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2238 VSS WL0[44] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2239 VSS WL0[44] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2240 VSS WL0[44] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2241 VSS WL0[44] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2242 VSS WL0[44] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2243 VSS WL0[44] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2244 VSS WL0[44] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2245 VSS WL0[44] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2246 VSS WL0[44] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2247 VSS WL0[44] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2248 VSS WL0[44] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2249 VSS WL0[44] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2250 VSS WL0[44] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2251 VSS WL0[44] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2252 VSS WL0[44] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2253 VSS WL0[44] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2254 VSS WL0[44] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2255 VSS WL0[44] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2256 VSS WL0[44] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2257 VSS WL0[44] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2258 VSS WL0[44] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2259 VSS WL0[44] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2260 VSS WL0[44] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2261 VSS WL0[44] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2262 VSS WL0[44] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2263 VSS WL0[44] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2264 VSS WL0[44] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2265 VSS WL0[44] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2266 VSS WL0[44] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2267 VSS WL0[44] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2268 VSS WL0[44] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2269 VSS WL0[44] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2270 VSS WL0[44] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2271 VSS WL0[44] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2272 VSS WL0[44] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2273 VSS WL0[44] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2274 VSS WL0[44] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2275 VSS WL0[44] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x2d0
XM2276 VSS WL0[45] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2277 VSS WL0[45] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2278 VSS WL0[45] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2279 VSS WL0[45] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2280 VSS WL0[45] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2281 VSS WL0[45] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2282 VSS WL0[45] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2283 VSS WL0[45] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2284 VSS WL0[45] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2285 VSS WL0[45] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2286 VSS WL0[45] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2287 VSS WL0[45] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2288 VSS WL0[45] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2289 VSS WL0[45] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2290 VSS WL0[45] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2291 VSS WL0[45] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2292 VSS WL0[45] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2293 VSS WL0[45] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2294 VSS WL0[45] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2295 VSS WL0[45] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2296 VSS WL0[45] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2297 VSS WL0[45] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2298 VSS WL0[45] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2299 VSS WL0[45] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2300 VSS WL0[45] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2301 VSS WL0[45] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2302 VSS WL0[45] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2303 VSS WL0[45] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2304 VSS WL0[45] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2305 VSS WL0[45] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2306 VSS WL0[45] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2307 VSS WL0[45] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2308 VSS WL0[45] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2309 VSS WL0[45] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2310 VSS WL0[45] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2311 VSS WL0[45] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2312 VSS WL0[45] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2313 VSS WL0[45] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2314 VSS WL0[45] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2315 VSS WL0[45] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2316 VSS WL0[45] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2317 VSS WL0[45] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2318 VSS WL0[45] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2319 VSS WL0[45] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2320 VSS WL0[45] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2321 VSS WL0[45] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2322 VSS WL0[45] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2323 VSS WL0[45] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2324 VSS WL0[45] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2325 VSS WL0[45] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2326 VSS WL0[45] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2327 VSS WL0[45] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2328 VSS WL0[45] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2329 VSS WL0[45] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2330 VSS WL0[45] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2331 VSS WL0[45] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2332 VSS WL0[45] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2333 VSS WL0[45] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2334 VSS WL0[45] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2335 VSS WL0[45] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2336 VSS WL0[45] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2337 VSS WL0[45] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2338 VSS WL0[45] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2339 VSS WL0[45] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2340 VSS WL0[45] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2341 VSS WL0[45] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2342 VSS WL0[45] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2343 VSS WL0[45] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x2e0
XM2344 VSS WL0[46] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2345 VSS WL0[46] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2346 VSS WL0[46] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2347 VSS WL0[46] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2348 VSS WL0[46] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2349 VSS WL0[46] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2350 VSS WL0[46] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2351 VSS WL0[46] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2352 VSS WL0[46] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2353 VSS WL0[46] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2354 VSS WL0[46] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2355 VSS WL0[46] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2356 VSS WL0[46] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2357 VSS WL0[46] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2358 VSS WL0[46] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2359 VSS WL0[46] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2360 VSS WL0[46] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2361 VSS WL0[46] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2362 VSS WL0[46] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2363 VSS WL0[46] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2364 VSS WL0[46] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2365 VSS WL0[46] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2366 VSS WL0[46] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2367 VSS WL0[46] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2368 VSS WL0[46] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2369 VSS WL0[46] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2370 VSS WL0[46] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2371 VSS WL0[46] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2372 VSS WL0[46] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2373 VSS WL0[46] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2374 VSS WL0[46] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2375 VSS WL0[46] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2376 VSS WL0[46] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2377 VSS WL0[46] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2378 VSS WL0[46] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2379 VSS WL0[46] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2380 VSS WL0[46] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2381 VSS WL0[46] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2382 VSS WL0[46] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2383 VSS WL0[46] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2384 VSS WL0[46] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2385 VSS WL0[46] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2386 VSS WL0[46] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2387 VSS WL0[46] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2388 VSS WL0[46] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2389 VSS WL0[46] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2390 VSS WL0[46] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2391 VSS WL0[46] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2392 VSS WL0[46] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2393 VSS WL0[46] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2394 VSS WL0[46] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2395 VSS WL0[46] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2396 VSS WL0[46] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2397 VSS WL0[46] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2398 VSS WL0[46] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2399 VSS WL0[46] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2400 VSS WL0[46] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2401 VSS WL0[46] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x2f0
XM2402 VSS WL0[47] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2403 VSS WL0[47] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2404 VSS WL0[47] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2405 VSS WL0[47] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2406 VSS WL0[47] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2407 VSS WL0[47] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2408 VSS WL0[47] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2409 VSS WL0[47] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2410 VSS WL0[47] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2411 VSS WL0[47] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2412 VSS WL0[47] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2413 VSS WL0[47] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2414 VSS WL0[47] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2415 VSS WL0[47] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2416 VSS WL0[47] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2417 VSS WL0[47] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2418 VSS WL0[47] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2419 VSS WL0[47] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2420 VSS WL0[47] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2421 VSS WL0[47] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2422 VSS WL0[47] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2423 VSS WL0[47] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2424 VSS WL0[47] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2425 VSS WL0[47] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2426 VSS WL0[47] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2427 VSS WL0[47] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2428 VSS WL0[47] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2429 VSS WL0[47] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2430 VSS WL0[47] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2431 VSS WL0[47] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2432 VSS WL0[47] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2433 VSS WL0[47] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2434 VSS WL0[47] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2435 VSS WL0[47] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2436 VSS WL0[47] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2437 VSS WL0[47] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2438 VSS WL0[47] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2439 VSS WL0[47] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2440 VSS WL0[47] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2441 VSS WL0[47] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2442 VSS WL0[47] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2443 VSS WL0[47] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2444 VSS WL0[47] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2445 VSS WL0[47] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2446 VSS WL0[47] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2447 VSS WL0[47] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2448 VSS WL0[47] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2449 VSS WL0[47] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x300
XM2450 VSS WL0[48] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2451 VSS WL0[48] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2452 VSS WL0[48] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2453 VSS WL0[48] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2454 VSS WL0[48] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2455 VSS WL0[48] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2456 VSS WL0[48] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2457 VSS WL0[48] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2458 VSS WL0[48] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2459 VSS WL0[48] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2460 VSS WL0[48] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2461 VSS WL0[48] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2462 VSS WL0[48] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2463 VSS WL0[48] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2464 VSS WL0[48] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2465 VSS WL0[48] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2466 VSS WL0[48] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2467 VSS WL0[48] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2468 VSS WL0[48] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2469 VSS WL0[48] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2470 VSS WL0[48] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2471 VSS WL0[48] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2472 VSS WL0[48] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2473 VSS WL0[48] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2474 VSS WL0[48] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2475 VSS WL0[48] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2476 VSS WL0[48] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2477 VSS WL0[48] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2478 VSS WL0[48] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2479 VSS WL0[48] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2480 VSS WL0[48] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2481 VSS WL0[48] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2482 VSS WL0[48] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2483 VSS WL0[48] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2484 VSS WL0[48] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2485 VSS WL0[48] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2486 VSS WL0[48] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2487 VSS WL0[48] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2488 VSS WL0[48] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2489 VSS WL0[48] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2490 VSS WL0[48] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2491 VSS WL0[48] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2492 VSS WL0[48] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2493 VSS WL0[48] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2494 VSS WL0[48] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2495 VSS WL0[48] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2496 VSS WL0[48] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2497 VSS WL0[48] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2498 VSS WL0[48] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2499 VSS WL0[48] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2500 VSS WL0[48] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x310
XM2501 VSS WL0[49] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2502 VSS WL0[49] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2503 VSS WL0[49] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2504 VSS WL0[49] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2505 VSS WL0[49] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2506 VSS WL0[49] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2507 VSS WL0[49] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2508 VSS WL0[49] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2509 VSS WL0[49] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2510 VSS WL0[49] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2511 VSS WL0[49] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2512 VSS WL0[49] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2513 VSS WL0[49] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2514 VSS WL0[49] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2515 VSS WL0[49] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2516 VSS WL0[49] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2517 VSS WL0[49] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2518 VSS WL0[49] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2519 VSS WL0[49] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2520 VSS WL0[49] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2521 VSS WL0[49] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2522 VSS WL0[49] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2523 VSS WL0[49] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2524 VSS WL0[49] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2525 VSS WL0[49] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2526 VSS WL0[49] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2527 VSS WL0[49] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2528 VSS WL0[49] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2529 VSS WL0[49] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2530 VSS WL0[49] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2531 VSS WL0[49] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2532 VSS WL0[49] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2533 VSS WL0[49] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2534 VSS WL0[49] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2535 VSS WL0[49] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2536 VSS WL0[49] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2537 VSS WL0[49] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2538 VSS WL0[49] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2539 VSS WL0[49] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2540 VSS WL0[49] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2541 VSS WL0[49] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2542 VSS WL0[49] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2543 VSS WL0[49] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2544 VSS WL0[49] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2545 VSS WL0[49] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2546 VSS WL0[49] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2547 VSS WL0[49] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2548 VSS WL0[49] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2549 VSS WL0[49] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2550 VSS WL0[49] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2551 VSS WL0[49] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2552 VSS WL0[49] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2553 VSS WL0[49] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2554 VSS WL0[49] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2555 VSS WL0[49] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2556 VSS WL0[49] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2557 VSS WL0[49] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2558 VSS WL0[49] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x320
XM2559 VSS WL0[50] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2560 VSS WL0[50] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2561 VSS WL0[50] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2562 VSS WL0[50] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2563 VSS WL0[50] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2564 VSS WL0[50] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2565 VSS WL0[50] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2566 VSS WL0[50] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2567 VSS WL0[50] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2568 VSS WL0[50] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2569 VSS WL0[50] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2570 VSS WL0[50] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2571 VSS WL0[50] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2572 VSS WL0[50] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2573 VSS WL0[50] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2574 VSS WL0[50] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2575 VSS WL0[50] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2576 VSS WL0[50] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2577 VSS WL0[50] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2578 VSS WL0[50] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2579 VSS WL0[50] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2580 VSS WL0[50] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2581 VSS WL0[50] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2582 VSS WL0[50] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2583 VSS WL0[50] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2584 VSS WL0[50] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2585 VSS WL0[50] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2586 VSS WL0[50] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2587 VSS WL0[50] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2588 VSS WL0[50] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2589 VSS WL0[50] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2590 VSS WL0[50] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2591 VSS WL0[50] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2592 VSS WL0[50] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2593 VSS WL0[50] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2594 VSS WL0[50] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2595 VSS WL0[50] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2596 VSS WL0[50] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2597 VSS WL0[50] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2598 VSS WL0[50] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2599 VSS WL0[50] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x330
XM2600 VSS WL0[51] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2601 VSS WL0[51] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2602 VSS WL0[51] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2603 VSS WL0[51] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2604 VSS WL0[51] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2605 VSS WL0[51] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2606 VSS WL0[51] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2607 VSS WL0[51] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2608 VSS WL0[51] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2609 VSS WL0[51] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2610 VSS WL0[51] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2611 VSS WL0[51] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2612 VSS WL0[51] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2613 VSS WL0[51] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2614 VSS WL0[51] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2615 VSS WL0[51] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2616 VSS WL0[51] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2617 VSS WL0[51] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2618 VSS WL0[51] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2619 VSS WL0[51] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2620 VSS WL0[51] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2621 VSS WL0[51] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2622 VSS WL0[51] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2623 VSS WL0[51] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2624 VSS WL0[51] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2625 VSS WL0[51] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2626 VSS WL0[51] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2627 VSS WL0[51] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2628 VSS WL0[51] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2629 VSS WL0[51] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2630 VSS WL0[51] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2631 VSS WL0[51] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2632 VSS WL0[51] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2633 VSS WL0[51] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2634 VSS WL0[51] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2635 VSS WL0[51] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2636 VSS WL0[51] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2637 VSS WL0[51] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2638 VSS WL0[51] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2639 VSS WL0[51] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2640 VSS WL0[51] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2641 VSS WL0[51] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2642 VSS WL0[51] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2643 VSS WL0[51] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2644 VSS WL0[51] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2645 VSS WL0[51] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2646 VSS WL0[51] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2647 VSS WL0[51] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2648 VSS WL0[51] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x340
XM2649 VSS WL0[52] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2650 VSS WL0[52] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2651 VSS WL0[52] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2652 VSS WL0[52] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2653 VSS WL0[52] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2654 VSS WL0[52] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2655 VSS WL0[52] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2656 VSS WL0[52] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2657 VSS WL0[52] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2658 VSS WL0[52] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2659 VSS WL0[52] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2660 VSS WL0[52] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2661 VSS WL0[52] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2662 VSS WL0[52] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2663 VSS WL0[52] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2664 VSS WL0[52] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2665 VSS WL0[52] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2666 VSS WL0[52] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2667 VSS WL0[52] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2668 VSS WL0[52] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2669 VSS WL0[52] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2670 VSS WL0[52] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2671 VSS WL0[52] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2672 VSS WL0[52] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2673 VSS WL0[52] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2674 VSS WL0[52] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2675 VSS WL0[52] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2676 VSS WL0[52] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2677 VSS WL0[52] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2678 VSS WL0[52] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2679 VSS WL0[52] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2680 VSS WL0[52] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2681 VSS WL0[52] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2682 VSS WL0[52] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2683 VSS WL0[52] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2684 VSS WL0[52] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2685 VSS WL0[52] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2686 VSS WL0[52] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2687 VSS WL0[52] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2688 VSS WL0[52] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2689 VSS WL0[52] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2690 VSS WL0[52] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2691 VSS WL0[52] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2692 VSS WL0[52] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2693 VSS WL0[52] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2694 VSS WL0[52] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2695 VSS WL0[52] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2696 VSS WL0[52] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2697 VSS WL0[52] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2698 VSS WL0[52] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2699 VSS WL0[52] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2700 VSS WL0[52] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2701 VSS WL0[52] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2702 VSS WL0[52] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2703 VSS WL0[52] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2704 VSS WL0[52] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2705 VSS WL0[52] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2706 VSS WL0[52] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2707 VSS WL0[52] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2708 VSS WL0[52] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2709 VSS WL0[52] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2710 VSS WL0[52] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2711 VSS WL0[52] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2712 VSS WL0[52] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2713 VSS WL0[52] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2714 VSS WL0[52] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x350
XM2715 VSS WL0[53] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2716 VSS WL0[53] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2717 VSS WL0[53] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2718 VSS WL0[53] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2719 VSS WL0[53] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2720 VSS WL0[53] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2721 VSS WL0[53] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2722 VSS WL0[53] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2723 VSS WL0[53] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2724 VSS WL0[53] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2725 VSS WL0[53] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2726 VSS WL0[53] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2727 VSS WL0[53] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2728 VSS WL0[53] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2729 VSS WL0[53] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2730 VSS WL0[53] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2731 VSS WL0[53] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2732 VSS WL0[53] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2733 VSS WL0[53] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2734 VSS WL0[53] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2735 VSS WL0[53] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2736 VSS WL0[53] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2737 VSS WL0[53] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2738 VSS WL0[53] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2739 VSS WL0[53] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2740 VSS WL0[53] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2741 VSS WL0[53] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2742 VSS WL0[53] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2743 VSS WL0[53] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2744 VSS WL0[53] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2745 VSS WL0[53] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2746 VSS WL0[53] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2747 VSS WL0[53] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2748 VSS WL0[53] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2749 VSS WL0[53] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2750 VSS WL0[53] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2751 VSS WL0[53] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2752 VSS WL0[53] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2753 VSS WL0[53] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2754 VSS WL0[53] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2755 VSS WL0[53] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2756 VSS WL0[53] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2757 VSS WL0[53] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2758 VSS WL0[53] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2759 VSS WL0[53] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2760 VSS WL0[53] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2761 VSS WL0[53] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2762 VSS WL0[53] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x360
XM2763 VSS WL0[54] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2764 VSS WL0[54] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2765 VSS WL0[54] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2766 VSS WL0[54] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2767 VSS WL0[54] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2768 VSS WL0[54] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2769 VSS WL0[54] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2770 VSS WL0[54] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2771 VSS WL0[54] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2772 VSS WL0[54] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2773 VSS WL0[54] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2774 VSS WL0[54] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2775 VSS WL0[54] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2776 VSS WL0[54] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2777 VSS WL0[54] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2778 VSS WL0[54] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2779 VSS WL0[54] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2780 VSS WL0[54] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2781 VSS WL0[54] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2782 VSS WL0[54] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2783 VSS WL0[54] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2784 VSS WL0[54] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2785 VSS WL0[54] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2786 VSS WL0[54] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2787 VSS WL0[54] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2788 VSS WL0[54] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2789 VSS WL0[54] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2790 VSS WL0[54] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2791 VSS WL0[54] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2792 VSS WL0[54] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2793 VSS WL0[54] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2794 VSS WL0[54] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2795 VSS WL0[54] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2796 VSS WL0[54] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2797 VSS WL0[54] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2798 VSS WL0[54] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2799 VSS WL0[54] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2800 VSS WL0[54] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2801 VSS WL0[54] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2802 VSS WL0[54] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2803 VSS WL0[54] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2804 VSS WL0[54] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2805 VSS WL0[54] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2806 VSS WL0[54] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2807 VSS WL0[54] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2808 VSS WL0[54] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2809 VSS WL0[54] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2810 VSS WL0[54] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2811 VSS WL0[54] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2812 VSS WL0[54] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2813 VSS WL0[54] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2814 VSS WL0[54] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2815 VSS WL0[54] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2816 VSS WL0[54] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2817 VSS WL0[54] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2818 VSS WL0[54] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2819 VSS WL0[54] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2820 VSS WL0[54] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2821 VSS WL0[54] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2822 VSS WL0[54] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2823 VSS WL0[54] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2824 VSS WL0[54] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2825 VSS WL0[54] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2826 VSS WL0[54] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2827 VSS WL0[54] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x370
XM2828 VSS WL0[55] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2829 VSS WL0[55] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2830 VSS WL0[55] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2831 VSS WL0[55] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2832 VSS WL0[55] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2833 VSS WL0[55] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2834 VSS WL0[55] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2835 VSS WL0[55] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2836 VSS WL0[55] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2837 VSS WL0[55] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2838 VSS WL0[55] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2839 VSS WL0[55] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2840 VSS WL0[55] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2841 VSS WL0[55] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2842 VSS WL0[55] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2843 VSS WL0[55] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2844 VSS WL0[55] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2845 VSS WL0[55] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2846 VSS WL0[55] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2847 VSS WL0[55] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2848 VSS WL0[55] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2849 VSS WL0[55] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2850 VSS WL0[55] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2851 VSS WL0[55] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2852 VSS WL0[55] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2853 VSS WL0[55] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2854 VSS WL0[55] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2855 VSS WL0[55] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2856 VSS WL0[55] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2857 VSS WL0[55] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2858 VSS WL0[55] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2859 VSS WL0[55] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2860 VSS WL0[55] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2861 VSS WL0[55] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2862 VSS WL0[55] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2863 VSS WL0[55] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2864 VSS WL0[55] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2865 VSS WL0[55] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2866 VSS WL0[55] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2867 VSS WL0[55] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2868 VSS WL0[55] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2869 VSS WL0[55] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2870 VSS WL0[55] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2871 VSS WL0[55] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2872 VSS WL0[55] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2873 VSS WL0[55] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2874 VSS WL0[55] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2875 VSS WL0[55] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2876 VSS WL0[55] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2877 VSS WL0[55] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2878 VSS WL0[55] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2879 VSS WL0[55] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2880 VSS WL0[55] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x380
XM2881 VSS WL0[56] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2882 VSS WL0[56] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2883 VSS WL0[56] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2884 VSS WL0[56] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2885 VSS WL0[56] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2886 VSS WL0[56] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2887 VSS WL0[56] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2888 VSS WL0[56] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2889 VSS WL0[56] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2890 VSS WL0[56] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2891 VSS WL0[56] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2892 VSS WL0[56] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2893 VSS WL0[56] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2894 VSS WL0[56] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2895 VSS WL0[56] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2896 VSS WL0[56] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2897 VSS WL0[56] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2898 VSS WL0[56] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2899 VSS WL0[56] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2900 VSS WL0[56] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2901 VSS WL0[56] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2902 VSS WL0[56] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2903 VSS WL0[56] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2904 VSS WL0[56] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2905 VSS WL0[56] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2906 VSS WL0[56] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2907 VSS WL0[56] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2908 VSS WL0[56] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2909 VSS WL0[56] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2910 VSS WL0[56] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2911 VSS WL0[56] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2912 VSS WL0[56] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2913 VSS WL0[56] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2914 VSS WL0[56] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2915 VSS WL0[56] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2916 VSS WL0[56] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2917 VSS WL0[56] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2918 VSS WL0[56] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2919 VSS WL0[56] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2920 VSS WL0[56] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2921 VSS WL0[56] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2922 VSS WL0[56] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2923 VSS WL0[56] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2924 VSS WL0[56] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2925 VSS WL0[56] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2926 VSS WL0[56] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2927 VSS WL0[56] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2928 VSS WL0[56] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2929 VSS WL0[56] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2930 VSS WL0[56] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2931 VSS WL0[56] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2932 VSS WL0[56] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2933 VSS WL0[56] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2934 VSS WL0[56] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2935 VSS WL0[56] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2936 VSS WL0[56] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x390
XM2937 VSS WL0[57] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2938 VSS WL0[57] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2939 VSS WL0[57] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2940 VSS WL0[57] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2941 VSS WL0[57] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2942 VSS WL0[57] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2943 VSS WL0[57] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2944 VSS WL0[57] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2945 VSS WL0[57] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2946 VSS WL0[57] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2947 VSS WL0[57] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2948 VSS WL0[57] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2949 VSS WL0[57] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2950 VSS WL0[57] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2951 VSS WL0[57] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2952 VSS WL0[57] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2953 VSS WL0[57] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2954 VSS WL0[57] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2955 VSS WL0[57] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2956 VSS WL0[57] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2957 VSS WL0[57] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2958 VSS WL0[57] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2959 VSS WL0[57] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2960 VSS WL0[57] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2961 VSS WL0[57] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2962 VSS WL0[57] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2963 VSS WL0[57] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2964 VSS WL0[57] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2965 VSS WL0[57] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2966 VSS WL0[57] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2967 VSS WL0[57] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2968 VSS WL0[57] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2969 VSS WL0[57] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2970 VSS WL0[57] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2971 VSS WL0[57] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2972 VSS WL0[57] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2973 VSS WL0[57] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2974 VSS WL0[57] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2975 VSS WL0[57] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2976 VSS WL0[57] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2977 VSS WL0[57] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2978 VSS WL0[57] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2979 VSS WL0[57] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2980 VSS WL0[57] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2981 VSS WL0[57] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2982 VSS WL0[57] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2983 VSS WL0[57] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2984 VSS WL0[57] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2985 VSS WL0[57] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2986 VSS WL0[57] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2987 VSS WL0[57] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2988 VSS WL0[57] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2989 VSS WL0[57] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2990 VSS WL0[57] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2991 VSS WL0[57] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2992 VSS WL0[57] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2993 VSS WL0[57] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2994 VSS WL0[57] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2995 VSS WL0[57] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2996 VSS WL0[57] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2997 VSS WL0[57] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM2998 VSS WL0[57] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x3a0
XM2999 VSS WL0[58] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3000 VSS WL0[58] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3001 VSS WL0[58] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3002 VSS WL0[58] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3003 VSS WL0[58] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3004 VSS WL0[58] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3005 VSS WL0[58] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3006 VSS WL0[58] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3007 VSS WL0[58] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3008 VSS WL0[58] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3009 VSS WL0[58] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3010 VSS WL0[58] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3011 VSS WL0[58] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3012 VSS WL0[58] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3013 VSS WL0[58] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3014 VSS WL0[58] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3015 VSS WL0[58] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3016 VSS WL0[58] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3017 VSS WL0[58] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3018 VSS WL0[58] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3019 VSS WL0[58] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3020 VSS WL0[58] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3021 VSS WL0[58] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3022 VSS WL0[58] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3023 VSS WL0[58] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3024 VSS WL0[58] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3025 VSS WL0[58] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3026 VSS WL0[58] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3027 VSS WL0[58] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3028 VSS WL0[58] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3029 VSS WL0[58] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3030 VSS WL0[58] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3031 VSS WL0[58] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3032 VSS WL0[58] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3033 VSS WL0[58] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3034 VSS WL0[58] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3035 VSS WL0[58] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3036 VSS WL0[58] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3037 VSS WL0[58] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3038 VSS WL0[58] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3039 VSS WL0[58] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3040 VSS WL0[58] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3041 VSS WL0[58] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3042 VSS WL0[58] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3043 VSS WL0[58] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3044 VSS WL0[58] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3045 VSS WL0[58] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3046 VSS WL0[58] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3047 VSS WL0[58] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3048 VSS WL0[58] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3049 VSS WL0[58] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3050 VSS WL0[58] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x3b0
XM3051 VSS WL0[59] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3052 VSS WL0[59] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3053 VSS WL0[59] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3054 VSS WL0[59] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3055 VSS WL0[59] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3056 VSS WL0[59] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3057 VSS WL0[59] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3058 VSS WL0[59] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3059 VSS WL0[59] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3060 VSS WL0[59] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3061 VSS WL0[59] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3062 VSS WL0[59] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3063 VSS WL0[59] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3064 VSS WL0[59] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3065 VSS WL0[59] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3066 VSS WL0[59] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3067 VSS WL0[59] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3068 VSS WL0[59] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3069 VSS WL0[59] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3070 VSS WL0[59] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3071 VSS WL0[59] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3072 VSS WL0[59] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3073 VSS WL0[59] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3074 VSS WL0[59] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3075 VSS WL0[59] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3076 VSS WL0[59] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3077 VSS WL0[59] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3078 VSS WL0[59] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3079 VSS WL0[59] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3080 VSS WL0[59] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3081 VSS WL0[59] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3082 VSS WL0[59] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3083 VSS WL0[59] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3084 VSS WL0[59] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3085 VSS WL0[59] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3086 VSS WL0[59] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3087 VSS WL0[59] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3088 VSS WL0[59] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3089 VSS WL0[59] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3090 VSS WL0[59] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3091 VSS WL0[59] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3092 VSS WL0[59] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3093 VSS WL0[59] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3094 VSS WL0[59] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3095 VSS WL0[59] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3096 VSS WL0[59] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3097 VSS WL0[59] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3098 VSS WL0[59] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3099 VSS WL0[59] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3100 VSS WL0[59] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3101 VSS WL0[59] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3102 VSS WL0[59] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3103 VSS WL0[59] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3104 VSS WL0[59] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3105 VSS WL0[59] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3106 VSS WL0[59] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3107 VSS WL0[59] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3108 VSS WL0[59] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3109 VSS WL0[59] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3110 VSS WL0[59] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3111 VSS WL0[59] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x3c0
XM3112 VSS WL0[60] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3113 VSS WL0[60] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3114 VSS WL0[60] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3115 VSS WL0[60] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3116 VSS WL0[60] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3117 VSS WL0[60] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3118 VSS WL0[60] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3119 VSS WL0[60] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3120 VSS WL0[60] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3121 VSS WL0[60] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3122 VSS WL0[60] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3123 VSS WL0[60] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3124 VSS WL0[60] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3125 VSS WL0[60] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3126 VSS WL0[60] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3127 VSS WL0[60] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3128 VSS WL0[60] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3129 VSS WL0[60] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3130 VSS WL0[60] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3131 VSS WL0[60] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3132 VSS WL0[60] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3133 VSS WL0[60] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3134 VSS WL0[60] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3135 VSS WL0[60] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3136 VSS WL0[60] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3137 VSS WL0[60] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3138 VSS WL0[60] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3139 VSS WL0[60] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3140 VSS WL0[60] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3141 VSS WL0[60] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3142 VSS WL0[60] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3143 VSS WL0[60] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3144 VSS WL0[60] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3145 VSS WL0[60] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3146 VSS WL0[60] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3147 VSS WL0[60] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3148 VSS WL0[60] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3149 VSS WL0[60] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3150 VSS WL0[60] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3151 VSS WL0[60] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3152 VSS WL0[60] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3153 VSS WL0[60] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3154 VSS WL0[60] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3155 VSS WL0[60] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3156 VSS WL0[60] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3157 VSS WL0[60] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3158 VSS WL0[60] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3159 VSS WL0[60] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3160 VSS WL0[60] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3161 VSS WL0[60] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3162 VSS WL0[60] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3163 VSS WL0[60] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3164 VSS WL0[60] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x3d0
XM3165 VSS WL0[61] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3166 VSS WL0[61] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3167 VSS WL0[61] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3168 VSS WL0[61] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3169 VSS WL0[61] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3170 VSS WL0[61] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3171 VSS WL0[61] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3172 VSS WL0[61] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3173 VSS WL0[61] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3174 VSS WL0[61] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3175 VSS WL0[61] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3176 VSS WL0[61] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3177 VSS WL0[61] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3178 VSS WL0[61] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3179 VSS WL0[61] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3180 VSS WL0[61] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3181 VSS WL0[61] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3182 VSS WL0[61] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3183 VSS WL0[61] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3184 VSS WL0[61] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3185 VSS WL0[61] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3186 VSS WL0[61] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3187 VSS WL0[61] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3188 VSS WL0[61] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3189 VSS WL0[61] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3190 VSS WL0[61] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3191 VSS WL0[61] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3192 VSS WL0[61] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3193 VSS WL0[61] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3194 VSS WL0[61] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3195 VSS WL0[61] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3196 VSS WL0[61] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3197 VSS WL0[61] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3198 VSS WL0[61] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3199 VSS WL0[61] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3200 VSS WL0[61] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3201 VSS WL0[61] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3202 VSS WL0[61] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3203 VSS WL0[61] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3204 VSS WL0[61] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3205 VSS WL0[61] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3206 VSS WL0[61] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3207 VSS WL0[61] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3208 VSS WL0[61] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3209 VSS WL0[61] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3210 VSS WL0[61] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3211 VSS WL0[61] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3212 VSS WL0[61] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3213 VSS WL0[61] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3214 VSS WL0[61] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3215 VSS WL0[61] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3216 VSS WL0[61] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3217 VSS WL0[61] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3218 VSS WL0[61] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3219 VSS WL0[61] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3220 VSS WL0[61] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3221 VSS WL0[61] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3222 VSS WL0[61] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3223 VSS WL0[61] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3224 VSS WL0[61] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3225 VSS WL0[61] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x3e0
XM3226 VSS WL0[62] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3227 VSS WL0[62] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3228 VSS WL0[62] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3229 VSS WL0[62] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3230 VSS WL0[62] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3231 VSS WL0[62] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3232 VSS WL0[62] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3233 VSS WL0[62] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3234 VSS WL0[62] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3235 VSS WL0[62] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3236 VSS WL0[62] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3237 VSS WL0[62] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3238 VSS WL0[62] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3239 VSS WL0[62] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3240 VSS WL0[62] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3241 VSS WL0[62] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3242 VSS WL0[62] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3243 VSS WL0[62] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3244 VSS WL0[62] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3245 VSS WL0[62] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3246 VSS WL0[62] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3247 VSS WL0[62] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3248 VSS WL0[62] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3249 VSS WL0[62] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3250 VSS WL0[62] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3251 VSS WL0[62] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3252 VSS WL0[62] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3253 VSS WL0[62] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3254 VSS WL0[62] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3255 VSS WL0[62] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3256 VSS WL0[62] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3257 VSS WL0[62] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3258 VSS WL0[62] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3259 VSS WL0[62] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3260 VSS WL0[62] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3261 VSS WL0[62] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3262 VSS WL0[62] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3263 VSS WL0[62] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3264 VSS WL0[62] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3265 VSS WL0[62] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3266 VSS WL0[62] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3267 VSS WL0[62] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3268 VSS WL0[62] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3269 VSS WL0[62] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3270 VSS WL0[62] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3271 VSS WL0[62] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3272 VSS WL0[62] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3273 VSS WL0[62] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3274 VSS WL0[62] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3275 VSS WL0[62] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x3f0
XM3276 VSS WL0[63] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3277 VSS WL0[63] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3278 VSS WL0[63] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3279 VSS WL0[63] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3280 VSS WL0[63] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3281 VSS WL0[63] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3282 VSS WL0[63] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3283 VSS WL0[63] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3284 VSS WL0[63] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3285 VSS WL0[63] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3286 VSS WL0[63] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3287 VSS WL0[63] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3288 VSS WL0[63] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3289 VSS WL0[63] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3290 VSS WL0[63] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3291 VSS WL0[63] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3292 VSS WL0[63] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3293 VSS WL0[63] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3294 VSS WL0[63] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3295 VSS WL0[63] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3296 VSS WL0[63] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3297 VSS WL0[63] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3298 VSS WL0[63] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3299 VSS WL0[63] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3300 VSS WL0[63] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3301 VSS WL0[63] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3302 VSS WL0[63] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3303 VSS WL0[63] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3304 VSS WL0[63] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3305 VSS WL0[63] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3306 VSS WL0[63] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3307 VSS WL0[63] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3308 VSS WL0[63] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3309 VSS WL0[63] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3310 VSS WL0[63] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3311 VSS WL0[63] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3312 VSS WL0[63] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3313 VSS WL0[63] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3314 VSS WL0[63] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3315 VSS WL0[63] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3316 VSS WL0[63] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3317 VSS WL0[63] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3318 VSS WL0[63] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3319 VSS WL0[63] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3320 VSS WL0[63] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3321 VSS WL0[63] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3322 VSS WL0[63] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3323 VSS WL0[63] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3324 VSS WL0[63] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3325 VSS WL0[63] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3326 VSS WL0[63] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3327 VSS WL0[63] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3328 VSS WL0[63] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3329 VSS WL0[63] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3330 VSS WL0[63] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3331 VSS WL0[63] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3332 VSS WL0[63] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3333 VSS WL0[63] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3334 VSS WL0[63] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3335 VSS WL0[63] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3336 VSS WL0[63] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3337 VSS WL0[63] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x400
XM3338 VSS WL0[64] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3339 VSS WL0[64] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3340 VSS WL0[64] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3341 VSS WL0[64] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3342 VSS WL0[64] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3343 VSS WL0[64] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3344 VSS WL0[64] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3345 VSS WL0[64] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3346 VSS WL0[64] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3347 VSS WL0[64] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3348 VSS WL0[64] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3349 VSS WL0[64] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3350 VSS WL0[64] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3351 VSS WL0[64] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3352 VSS WL0[64] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3353 VSS WL0[64] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3354 VSS WL0[64] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3355 VSS WL0[64] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3356 VSS WL0[64] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3357 VSS WL0[64] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3358 VSS WL0[64] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3359 VSS WL0[64] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3360 VSS WL0[64] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3361 VSS WL0[64] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3362 VSS WL0[64] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3363 VSS WL0[64] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3364 VSS WL0[64] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3365 VSS WL0[64] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3366 VSS WL0[64] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3367 VSS WL0[64] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3368 VSS WL0[64] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3369 VSS WL0[64] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3370 VSS WL0[64] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3371 VSS WL0[64] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3372 VSS WL0[64] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3373 VSS WL0[64] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3374 VSS WL0[64] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3375 VSS WL0[64] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3376 VSS WL0[64] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3377 VSS WL0[64] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3378 VSS WL0[64] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3379 VSS WL0[64] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3380 VSS WL0[64] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3381 VSS WL0[64] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3382 VSS WL0[64] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3383 VSS WL0[64] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3384 VSS WL0[64] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3385 VSS WL0[64] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3386 VSS WL0[64] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3387 VSS WL0[64] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3388 VSS WL0[64] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3389 VSS WL0[64] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3390 VSS WL0[64] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3391 VSS WL0[64] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x410
XM3392 VSS WL0[65] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3393 VSS WL0[65] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3394 VSS WL0[65] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3395 VSS WL0[65] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3396 VSS WL0[65] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3397 VSS WL0[65] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3398 VSS WL0[65] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3399 VSS WL0[65] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3400 VSS WL0[65] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3401 VSS WL0[65] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3402 VSS WL0[65] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3403 VSS WL0[65] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3404 VSS WL0[65] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3405 VSS WL0[65] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3406 VSS WL0[65] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3407 VSS WL0[65] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3408 VSS WL0[65] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3409 VSS WL0[65] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3410 VSS WL0[65] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3411 VSS WL0[65] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3412 VSS WL0[65] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3413 VSS WL0[65] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3414 VSS WL0[65] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3415 VSS WL0[65] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3416 VSS WL0[65] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3417 VSS WL0[65] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3418 VSS WL0[65] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3419 VSS WL0[65] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3420 VSS WL0[65] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3421 VSS WL0[65] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3422 VSS WL0[65] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3423 VSS WL0[65] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3424 VSS WL0[65] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3425 VSS WL0[65] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3426 VSS WL0[65] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3427 VSS WL0[65] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3428 VSS WL0[65] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3429 VSS WL0[65] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3430 VSS WL0[65] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3431 VSS WL0[65] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3432 VSS WL0[65] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3433 VSS WL0[65] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3434 VSS WL0[65] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3435 VSS WL0[65] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3436 VSS WL0[65] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3437 VSS WL0[65] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3438 VSS WL0[65] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3439 VSS WL0[65] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3440 VSS WL0[65] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3441 VSS WL0[65] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3442 VSS WL0[65] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3443 VSS WL0[65] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3444 VSS WL0[65] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3445 VSS WL0[65] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x420
XM3446 VSS WL0[66] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3447 VSS WL0[66] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3448 VSS WL0[66] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3449 VSS WL0[66] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3450 VSS WL0[66] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3451 VSS WL0[66] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3452 VSS WL0[66] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3453 VSS WL0[66] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3454 VSS WL0[66] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3455 VSS WL0[66] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3456 VSS WL0[66] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3457 VSS WL0[66] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3458 VSS WL0[66] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3459 VSS WL0[66] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3460 VSS WL0[66] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3461 VSS WL0[66] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3462 VSS WL0[66] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3463 VSS WL0[66] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3464 VSS WL0[66] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3465 VSS WL0[66] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3466 VSS WL0[66] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3467 VSS WL0[66] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3468 VSS WL0[66] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3469 VSS WL0[66] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3470 VSS WL0[66] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3471 VSS WL0[66] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3472 VSS WL0[66] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3473 VSS WL0[66] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3474 VSS WL0[66] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3475 VSS WL0[66] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3476 VSS WL0[66] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3477 VSS WL0[66] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3478 VSS WL0[66] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3479 VSS WL0[66] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3480 VSS WL0[66] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3481 VSS WL0[66] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3482 VSS WL0[66] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3483 VSS WL0[66] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3484 VSS WL0[66] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3485 VSS WL0[66] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3486 VSS WL0[66] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3487 VSS WL0[66] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3488 VSS WL0[66] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3489 VSS WL0[66] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3490 VSS WL0[66] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3491 VSS WL0[66] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3492 VSS WL0[66] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3493 VSS WL0[66] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3494 VSS WL0[66] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3495 VSS WL0[66] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3496 VSS WL0[66] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3497 VSS WL0[66] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3498 VSS WL0[66] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3499 VSS WL0[66] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3500 VSS WL0[66] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3501 VSS WL0[66] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3502 VSS WL0[66] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3503 VSS WL0[66] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3504 VSS WL0[66] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3505 VSS WL0[66] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3506 VSS WL0[66] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3507 VSS WL0[66] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x430
XM3508 VSS WL0[67] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3509 VSS WL0[67] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3510 VSS WL0[67] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3511 VSS WL0[67] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3512 VSS WL0[67] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3513 VSS WL0[67] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3514 VSS WL0[67] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3515 VSS WL0[67] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3516 VSS WL0[67] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3517 VSS WL0[67] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3518 VSS WL0[67] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3519 VSS WL0[67] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3520 VSS WL0[67] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3521 VSS WL0[67] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3522 VSS WL0[67] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3523 VSS WL0[67] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3524 VSS WL0[67] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3525 VSS WL0[67] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3526 VSS WL0[67] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3527 VSS WL0[67] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3528 VSS WL0[67] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3529 VSS WL0[67] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3530 VSS WL0[67] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3531 VSS WL0[67] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3532 VSS WL0[67] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3533 VSS WL0[67] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3534 VSS WL0[67] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3535 VSS WL0[67] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3536 VSS WL0[67] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3537 VSS WL0[67] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3538 VSS WL0[67] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3539 VSS WL0[67] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3540 VSS WL0[67] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3541 VSS WL0[67] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3542 VSS WL0[67] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3543 VSS WL0[67] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3544 VSS WL0[67] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3545 VSS WL0[67] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3546 VSS WL0[67] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3547 VSS WL0[67] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3548 VSS WL0[67] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3549 VSS WL0[67] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3550 VSS WL0[67] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3551 VSS WL0[67] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3552 VSS WL0[67] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3553 VSS WL0[67] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3554 VSS WL0[67] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3555 VSS WL0[67] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3556 VSS WL0[67] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3557 VSS WL0[67] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3558 VSS WL0[67] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x440
XM3559 VSS WL0[68] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3560 VSS WL0[68] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3561 VSS WL0[68] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3562 VSS WL0[68] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3563 VSS WL0[68] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3564 VSS WL0[68] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3565 VSS WL0[68] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3566 VSS WL0[68] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3567 VSS WL0[68] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3568 VSS WL0[68] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3569 VSS WL0[68] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3570 VSS WL0[68] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3571 VSS WL0[68] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3572 VSS WL0[68] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3573 VSS WL0[68] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3574 VSS WL0[68] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3575 VSS WL0[68] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3576 VSS WL0[68] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3577 VSS WL0[68] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3578 VSS WL0[68] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3579 VSS WL0[68] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3580 VSS WL0[68] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3581 VSS WL0[68] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3582 VSS WL0[68] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3583 VSS WL0[68] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3584 VSS WL0[68] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3585 VSS WL0[68] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3586 VSS WL0[68] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3587 VSS WL0[68] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3588 VSS WL0[68] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3589 VSS WL0[68] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3590 VSS WL0[68] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3591 VSS WL0[68] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3592 VSS WL0[68] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3593 VSS WL0[68] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3594 VSS WL0[68] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3595 VSS WL0[68] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3596 VSS WL0[68] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3597 VSS WL0[68] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3598 VSS WL0[68] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3599 VSS WL0[68] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3600 VSS WL0[68] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3601 VSS WL0[68] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3602 VSS WL0[68] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3603 VSS WL0[68] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3604 VSS WL0[68] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3605 VSS WL0[68] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3606 VSS WL0[68] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3607 VSS WL0[68] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3608 VSS WL0[68] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3609 VSS WL0[68] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3610 VSS WL0[68] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3611 VSS WL0[68] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3612 VSS WL0[68] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3613 VSS WL0[68] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3614 VSS WL0[68] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3615 VSS WL0[68] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3616 VSS WL0[68] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3617 VSS WL0[68] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3618 VSS WL0[68] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3619 VSS WL0[68] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x450
XM3620 VSS WL0[69] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3621 VSS WL0[69] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3622 VSS WL0[69] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3623 VSS WL0[69] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3624 VSS WL0[69] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3625 VSS WL0[69] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3626 VSS WL0[69] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3627 VSS WL0[69] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3628 VSS WL0[69] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3629 VSS WL0[69] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3630 VSS WL0[69] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3631 VSS WL0[69] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3632 VSS WL0[69] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3633 VSS WL0[69] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3634 VSS WL0[69] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3635 VSS WL0[69] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3636 VSS WL0[69] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3637 VSS WL0[69] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3638 VSS WL0[69] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3639 VSS WL0[69] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3640 VSS WL0[69] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3641 VSS WL0[69] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3642 VSS WL0[69] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3643 VSS WL0[69] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3644 VSS WL0[69] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3645 VSS WL0[69] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3646 VSS WL0[69] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3647 VSS WL0[69] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3648 VSS WL0[69] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3649 VSS WL0[69] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3650 VSS WL0[69] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3651 VSS WL0[69] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3652 VSS WL0[69] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3653 VSS WL0[69] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3654 VSS WL0[69] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3655 VSS WL0[69] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3656 VSS WL0[69] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3657 VSS WL0[69] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3658 VSS WL0[69] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3659 VSS WL0[69] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3660 VSS WL0[69] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3661 VSS WL0[69] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3662 VSS WL0[69] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3663 VSS WL0[69] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3664 VSS WL0[69] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3665 VSS WL0[69] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3666 VSS WL0[69] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3667 VSS WL0[69] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3668 VSS WL0[69] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3669 VSS WL0[69] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3670 VSS WL0[69] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x460
XM3671 VSS WL0[70] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3672 VSS WL0[70] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3673 VSS WL0[70] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3674 VSS WL0[70] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3675 VSS WL0[70] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3676 VSS WL0[70] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3677 VSS WL0[70] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3678 VSS WL0[70] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3679 VSS WL0[70] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3680 VSS WL0[70] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3681 VSS WL0[70] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3682 VSS WL0[70] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3683 VSS WL0[70] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3684 VSS WL0[70] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3685 VSS WL0[70] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3686 VSS WL0[70] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3687 VSS WL0[70] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3688 VSS WL0[70] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3689 VSS WL0[70] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3690 VSS WL0[70] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3691 VSS WL0[70] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3692 VSS WL0[70] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3693 VSS WL0[70] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3694 VSS WL0[70] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3695 VSS WL0[70] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3696 VSS WL0[70] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3697 VSS WL0[70] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3698 VSS WL0[70] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3699 VSS WL0[70] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3700 VSS WL0[70] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3701 VSS WL0[70] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3702 VSS WL0[70] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3703 VSS WL0[70] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3704 VSS WL0[70] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3705 VSS WL0[70] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3706 VSS WL0[70] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3707 VSS WL0[70] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3708 VSS WL0[70] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3709 VSS WL0[70] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3710 VSS WL0[70] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3711 VSS WL0[70] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3712 VSS WL0[70] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3713 VSS WL0[70] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3714 VSS WL0[70] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3715 VSS WL0[70] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3716 VSS WL0[70] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3717 VSS WL0[70] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3718 VSS WL0[70] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3719 VSS WL0[70] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3720 VSS WL0[70] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3721 VSS WL0[70] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3722 VSS WL0[70] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3723 VSS WL0[70] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3724 VSS WL0[70] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3725 VSS WL0[70] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3726 VSS WL0[70] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3727 VSS WL0[70] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3728 VSS WL0[70] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3729 VSS WL0[70] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3730 VSS WL0[70] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3731 VSS WL0[70] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x470
XM3732 VSS WL0[71] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3733 VSS WL0[71] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3734 VSS WL0[71] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3735 VSS WL0[71] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3736 VSS WL0[71] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3737 VSS WL0[71] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3738 VSS WL0[71] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3739 VSS WL0[71] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3740 VSS WL0[71] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3741 VSS WL0[71] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3742 VSS WL0[71] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3743 VSS WL0[71] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3744 VSS WL0[71] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3745 VSS WL0[71] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3746 VSS WL0[71] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3747 VSS WL0[71] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3748 VSS WL0[71] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3749 VSS WL0[71] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3750 VSS WL0[71] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3751 VSS WL0[71] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3752 VSS WL0[71] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3753 VSS WL0[71] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3754 VSS WL0[71] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3755 VSS WL0[71] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3756 VSS WL0[71] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3757 VSS WL0[71] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3758 VSS WL0[71] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3759 VSS WL0[71] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3760 VSS WL0[71] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3761 VSS WL0[71] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3762 VSS WL0[71] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3763 VSS WL0[71] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3764 VSS WL0[71] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3765 VSS WL0[71] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3766 VSS WL0[71] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3767 VSS WL0[71] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3768 VSS WL0[71] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3769 VSS WL0[71] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3770 VSS WL0[71] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3771 VSS WL0[71] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3772 VSS WL0[71] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3773 VSS WL0[71] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3774 VSS WL0[71] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3775 VSS WL0[71] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3776 VSS WL0[71] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3777 VSS WL0[71] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3778 VSS WL0[71] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3779 VSS WL0[71] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3780 VSS WL0[71] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3781 VSS WL0[71] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3782 VSS WL0[71] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x480
XM3783 VSS WL0[72] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3784 VSS WL0[72] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3785 VSS WL0[72] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3786 VSS WL0[72] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3787 VSS WL0[72] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3788 VSS WL0[72] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3789 VSS WL0[72] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3790 VSS WL0[72] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3791 VSS WL0[72] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3792 VSS WL0[72] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3793 VSS WL0[72] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3794 VSS WL0[72] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3795 VSS WL0[72] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3796 VSS WL0[72] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3797 VSS WL0[72] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3798 VSS WL0[72] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3799 VSS WL0[72] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3800 VSS WL0[72] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3801 VSS WL0[72] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3802 VSS WL0[72] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3803 VSS WL0[72] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3804 VSS WL0[72] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3805 VSS WL0[72] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3806 VSS WL0[72] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3807 VSS WL0[72] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3808 VSS WL0[72] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3809 VSS WL0[72] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3810 VSS WL0[72] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3811 VSS WL0[72] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3812 VSS WL0[72] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3813 VSS WL0[72] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3814 VSS WL0[72] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3815 VSS WL0[72] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3816 VSS WL0[72] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3817 VSS WL0[72] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3818 VSS WL0[72] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3819 VSS WL0[72] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3820 VSS WL0[72] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3821 VSS WL0[72] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3822 VSS WL0[72] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3823 VSS WL0[72] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3824 VSS WL0[72] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3825 VSS WL0[72] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3826 VSS WL0[72] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3827 VSS WL0[72] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3828 VSS WL0[72] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3829 VSS WL0[72] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3830 VSS WL0[72] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3831 VSS WL0[72] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3832 VSS WL0[72] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3833 VSS WL0[72] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3834 VSS WL0[72] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3835 VSS WL0[72] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3836 VSS WL0[72] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3837 VSS WL0[72] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3838 VSS WL0[72] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3839 VSS WL0[72] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3840 VSS WL0[72] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3841 VSS WL0[72] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3842 VSS WL0[72] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3843 VSS WL0[72] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x490
XM3844 VSS WL0[73] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3845 VSS WL0[73] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3846 VSS WL0[73] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3847 VSS WL0[73] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3848 VSS WL0[73] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3849 VSS WL0[73] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3850 VSS WL0[73] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3851 VSS WL0[73] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3852 VSS WL0[73] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3853 VSS WL0[73] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3854 VSS WL0[73] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3855 VSS WL0[73] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3856 VSS WL0[73] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3857 VSS WL0[73] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3858 VSS WL0[73] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3859 VSS WL0[73] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3860 VSS WL0[73] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3861 VSS WL0[73] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3862 VSS WL0[73] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3863 VSS WL0[73] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3864 VSS WL0[73] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3865 VSS WL0[73] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3866 VSS WL0[73] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3867 VSS WL0[73] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3868 VSS WL0[73] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3869 VSS WL0[73] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3870 VSS WL0[73] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3871 VSS WL0[73] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3872 VSS WL0[73] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3873 VSS WL0[73] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3874 VSS WL0[73] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3875 VSS WL0[73] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3876 VSS WL0[73] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3877 VSS WL0[73] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3878 VSS WL0[73] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3879 VSS WL0[73] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3880 VSS WL0[73] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3881 VSS WL0[73] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3882 VSS WL0[73] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3883 VSS WL0[73] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3884 VSS WL0[73] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3885 VSS WL0[73] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3886 VSS WL0[73] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3887 VSS WL0[73] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3888 VSS WL0[73] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3889 VSS WL0[73] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3890 VSS WL0[73] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3891 VSS WL0[73] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3892 VSS WL0[73] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3893 VSS WL0[73] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3894 VSS WL0[73] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3895 VSS WL0[73] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3896 VSS WL0[73] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3897 VSS WL0[73] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x4a0
XM3898 VSS WL0[74] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3899 VSS WL0[74] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3900 VSS WL0[74] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3901 VSS WL0[74] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3902 VSS WL0[74] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3903 VSS WL0[74] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3904 VSS WL0[74] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3905 VSS WL0[74] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3906 VSS WL0[74] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3907 VSS WL0[74] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3908 VSS WL0[74] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3909 VSS WL0[74] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3910 VSS WL0[74] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3911 VSS WL0[74] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3912 VSS WL0[74] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3913 VSS WL0[74] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3914 VSS WL0[74] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3915 VSS WL0[74] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3916 VSS WL0[74] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3917 VSS WL0[74] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3918 VSS WL0[74] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3919 VSS WL0[74] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3920 VSS WL0[74] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3921 VSS WL0[74] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3922 VSS WL0[74] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3923 VSS WL0[74] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3924 VSS WL0[74] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3925 VSS WL0[74] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3926 VSS WL0[74] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3927 VSS WL0[74] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3928 VSS WL0[74] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3929 VSS WL0[74] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3930 VSS WL0[74] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3931 VSS WL0[74] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3932 VSS WL0[74] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3933 VSS WL0[74] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3934 VSS WL0[74] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3935 VSS WL0[74] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3936 VSS WL0[74] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3937 VSS WL0[74] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3938 VSS WL0[74] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3939 VSS WL0[74] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3940 VSS WL0[74] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3941 VSS WL0[74] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3942 VSS WL0[74] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3943 VSS WL0[74] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3944 VSS WL0[74] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3945 VSS WL0[74] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3946 VSS WL0[74] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3947 VSS WL0[74] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3948 VSS WL0[74] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3949 VSS WL0[74] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3950 VSS WL0[74] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3951 VSS WL0[74] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x4b0
XM3952 VSS WL0[75] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3953 VSS WL0[75] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3954 VSS WL0[75] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3955 VSS WL0[75] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3956 VSS WL0[75] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3957 VSS WL0[75] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3958 VSS WL0[75] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3959 VSS WL0[75] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3960 VSS WL0[75] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3961 VSS WL0[75] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3962 VSS WL0[75] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3963 VSS WL0[75] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3964 VSS WL0[75] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3965 VSS WL0[75] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3966 VSS WL0[75] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3967 VSS WL0[75] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3968 VSS WL0[75] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3969 VSS WL0[75] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3970 VSS WL0[75] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3971 VSS WL0[75] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3972 VSS WL0[75] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3973 VSS WL0[75] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3974 VSS WL0[75] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3975 VSS WL0[75] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3976 VSS WL0[75] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3977 VSS WL0[75] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3978 VSS WL0[75] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3979 VSS WL0[75] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3980 VSS WL0[75] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3981 VSS WL0[75] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3982 VSS WL0[75] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3983 VSS WL0[75] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3984 VSS WL0[75] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3985 VSS WL0[75] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3986 VSS WL0[75] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3987 VSS WL0[75] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3988 VSS WL0[75] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3989 VSS WL0[75] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3990 VSS WL0[75] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3991 VSS WL0[75] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3992 VSS WL0[75] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3993 VSS WL0[75] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3994 VSS WL0[75] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3995 VSS WL0[75] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3996 VSS WL0[75] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3997 VSS WL0[75] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3998 VSS WL0[75] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM3999 VSS WL0[75] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4000 VSS WL0[75] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4001 VSS WL0[75] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4002 VSS WL0[75] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4003 VSS WL0[75] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4004 VSS WL0[75] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4005 VSS WL0[75] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4006 VSS WL0[75] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4007 VSS WL0[75] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4008 VSS WL0[75] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4009 VSS WL0[75] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4010 VSS WL0[75] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4011 VSS WL0[75] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4012 VSS WL0[75] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4013 VSS WL0[75] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x4c0
XM4014 VSS WL0[76] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4015 VSS WL0[76] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4016 VSS WL0[76] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4017 VSS WL0[76] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4018 VSS WL0[76] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4019 VSS WL0[76] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4020 VSS WL0[76] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4021 VSS WL0[76] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4022 VSS WL0[76] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4023 VSS WL0[76] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4024 VSS WL0[76] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4025 VSS WL0[76] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4026 VSS WL0[76] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4027 VSS WL0[76] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4028 VSS WL0[76] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4029 VSS WL0[76] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4030 VSS WL0[76] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4031 VSS WL0[76] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4032 VSS WL0[76] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4033 VSS WL0[76] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4034 VSS WL0[76] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4035 VSS WL0[76] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4036 VSS WL0[76] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4037 VSS WL0[76] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4038 VSS WL0[76] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4039 VSS WL0[76] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4040 VSS WL0[76] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4041 VSS WL0[76] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4042 VSS WL0[76] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4043 VSS WL0[76] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4044 VSS WL0[76] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4045 VSS WL0[76] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4046 VSS WL0[76] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4047 VSS WL0[76] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4048 VSS WL0[76] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4049 VSS WL0[76] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4050 VSS WL0[76] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4051 VSS WL0[76] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4052 VSS WL0[76] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4053 VSS WL0[76] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4054 VSS WL0[76] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4055 VSS WL0[76] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4056 VSS WL0[76] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4057 VSS WL0[76] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4058 VSS WL0[76] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4059 VSS WL0[76] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4060 VSS WL0[76] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4061 VSS WL0[76] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4062 VSS WL0[76] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4063 VSS WL0[76] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4064 VSS WL0[76] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4065 VSS WL0[76] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x4d0
XM4066 VSS WL0[77] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4067 VSS WL0[77] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4068 VSS WL0[77] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4069 VSS WL0[77] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4070 VSS WL0[77] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4071 VSS WL0[77] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4072 VSS WL0[77] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4073 VSS WL0[77] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4074 VSS WL0[77] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4075 VSS WL0[77] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4076 VSS WL0[77] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4077 VSS WL0[77] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4078 VSS WL0[77] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4079 VSS WL0[77] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4080 VSS WL0[77] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4081 VSS WL0[77] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4082 VSS WL0[77] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4083 VSS WL0[77] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4084 VSS WL0[77] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4085 VSS WL0[77] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4086 VSS WL0[77] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4087 VSS WL0[77] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4088 VSS WL0[77] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4089 VSS WL0[77] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4090 VSS WL0[77] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4091 VSS WL0[77] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4092 VSS WL0[77] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4093 VSS WL0[77] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4094 VSS WL0[77] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4095 VSS WL0[77] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4096 VSS WL0[77] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4097 VSS WL0[77] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4098 VSS WL0[77] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4099 VSS WL0[77] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4100 VSS WL0[77] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4101 VSS WL0[77] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4102 VSS WL0[77] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4103 VSS WL0[77] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4104 VSS WL0[77] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4105 VSS WL0[77] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4106 VSS WL0[77] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4107 VSS WL0[77] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4108 VSS WL0[77] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4109 VSS WL0[77] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4110 VSS WL0[77] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4111 VSS WL0[77] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4112 VSS WL0[77] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4113 VSS WL0[77] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4114 VSS WL0[77] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4115 VSS WL0[77] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4116 VSS WL0[77] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4117 VSS WL0[77] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4118 VSS WL0[77] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4119 VSS WL0[77] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4120 VSS WL0[77] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4121 VSS WL0[77] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4122 VSS WL0[77] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4123 VSS WL0[77] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4124 VSS WL0[77] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4125 VSS WL0[77] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4126 VSS WL0[77] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x4e0
XM4127 VSS WL0[78] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4128 VSS WL0[78] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4129 VSS WL0[78] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4130 VSS WL0[78] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4131 VSS WL0[78] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4132 VSS WL0[78] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4133 VSS WL0[78] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4134 VSS WL0[78] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4135 VSS WL0[78] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4136 VSS WL0[78] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4137 VSS WL0[78] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4138 VSS WL0[78] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4139 VSS WL0[78] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4140 VSS WL0[78] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4141 VSS WL0[78] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4142 VSS WL0[78] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4143 VSS WL0[78] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4144 VSS WL0[78] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4145 VSS WL0[78] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4146 VSS WL0[78] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4147 VSS WL0[78] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4148 VSS WL0[78] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4149 VSS WL0[78] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4150 VSS WL0[78] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4151 VSS WL0[78] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4152 VSS WL0[78] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4153 VSS WL0[78] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4154 VSS WL0[78] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4155 VSS WL0[78] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4156 VSS WL0[78] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4157 VSS WL0[78] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4158 VSS WL0[78] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4159 VSS WL0[78] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4160 VSS WL0[78] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4161 VSS WL0[78] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4162 VSS WL0[78] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4163 VSS WL0[78] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4164 VSS WL0[78] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4165 VSS WL0[78] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4166 VSS WL0[78] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4167 VSS WL0[78] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4168 VSS WL0[78] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4169 VSS WL0[78] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4170 VSS WL0[78] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4171 VSS WL0[78] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4172 VSS WL0[78] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4173 VSS WL0[78] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4174 VSS WL0[78] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4175 VSS WL0[78] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4176 VSS WL0[78] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4177 VSS WL0[78] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4178 VSS WL0[78] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x4f0
XM4179 VSS WL0[79] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4180 VSS WL0[79] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4181 VSS WL0[79] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4182 VSS WL0[79] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4183 VSS WL0[79] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4184 VSS WL0[79] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4185 VSS WL0[79] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4186 VSS WL0[79] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4187 VSS WL0[79] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4188 VSS WL0[79] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4189 VSS WL0[79] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4190 VSS WL0[79] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4191 VSS WL0[79] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4192 VSS WL0[79] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4193 VSS WL0[79] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4194 VSS WL0[79] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4195 VSS WL0[79] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4196 VSS WL0[79] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4197 VSS WL0[79] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4198 VSS WL0[79] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4199 VSS WL0[79] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4200 VSS WL0[79] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4201 VSS WL0[79] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4202 VSS WL0[79] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4203 VSS WL0[79] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4204 VSS WL0[79] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4205 VSS WL0[79] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4206 VSS WL0[79] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4207 VSS WL0[79] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4208 VSS WL0[79] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4209 VSS WL0[79] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4210 VSS WL0[79] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4211 VSS WL0[79] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4212 VSS WL0[79] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4213 VSS WL0[79] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4214 VSS WL0[79] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4215 VSS WL0[79] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4216 VSS WL0[79] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4217 VSS WL0[79] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4218 VSS WL0[79] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4219 VSS WL0[79] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4220 VSS WL0[79] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4221 VSS WL0[79] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4222 VSS WL0[79] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4223 VSS WL0[79] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4224 VSS WL0[79] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4225 VSS WL0[79] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4226 VSS WL0[79] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4227 VSS WL0[79] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4228 VSS WL0[79] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4229 VSS WL0[79] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4230 VSS WL0[79] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4231 VSS WL0[79] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4232 VSS WL0[79] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4233 VSS WL0[79] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4234 VSS WL0[79] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4235 VSS WL0[79] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4236 VSS WL0[79] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4237 VSS WL0[79] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4238 VSS WL0[79] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4239 VSS WL0[79] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x500
XM4240 VSS WL0[80] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4241 VSS WL0[80] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4242 VSS WL0[80] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4243 VSS WL0[80] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4244 VSS WL0[80] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4245 VSS WL0[80] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4246 VSS WL0[80] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4247 VSS WL0[80] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4248 VSS WL0[80] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4249 VSS WL0[80] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4250 VSS WL0[80] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4251 VSS WL0[80] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4252 VSS WL0[80] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4253 VSS WL0[80] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4254 VSS WL0[80] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4255 VSS WL0[80] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4256 VSS WL0[80] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4257 VSS WL0[80] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4258 VSS WL0[80] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4259 VSS WL0[80] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4260 VSS WL0[80] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4261 VSS WL0[80] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4262 VSS WL0[80] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4263 VSS WL0[80] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4264 VSS WL0[80] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4265 VSS WL0[80] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4266 VSS WL0[80] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4267 VSS WL0[80] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4268 VSS WL0[80] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4269 VSS WL0[80] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4270 VSS WL0[80] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4271 VSS WL0[80] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4272 VSS WL0[80] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4273 VSS WL0[80] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4274 VSS WL0[80] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4275 VSS WL0[80] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4276 VSS WL0[80] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4277 VSS WL0[80] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4278 VSS WL0[80] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4279 VSS WL0[80] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4280 VSS WL0[80] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4281 VSS WL0[80] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4282 VSS WL0[80] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4283 VSS WL0[80] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4284 VSS WL0[80] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4285 VSS WL0[80] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4286 VSS WL0[80] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4287 VSS WL0[80] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4288 VSS WL0[80] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4289 VSS WL0[80] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4290 VSS WL0[80] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4291 VSS WL0[80] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x510
XM4292 VSS WL0[81] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4293 VSS WL0[81] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4294 VSS WL0[81] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4295 VSS WL0[81] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4296 VSS WL0[81] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4297 VSS WL0[81] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4298 VSS WL0[81] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4299 VSS WL0[81] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4300 VSS WL0[81] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4301 VSS WL0[81] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4302 VSS WL0[81] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4303 VSS WL0[81] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4304 VSS WL0[81] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4305 VSS WL0[81] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4306 VSS WL0[81] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4307 VSS WL0[81] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4308 VSS WL0[81] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4309 VSS WL0[81] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4310 VSS WL0[81] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4311 VSS WL0[81] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4312 VSS WL0[81] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4313 VSS WL0[81] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4314 VSS WL0[81] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4315 VSS WL0[81] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4316 VSS WL0[81] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4317 VSS WL0[81] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4318 VSS WL0[81] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4319 VSS WL0[81] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4320 VSS WL0[81] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4321 VSS WL0[81] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4322 VSS WL0[81] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4323 VSS WL0[81] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4324 VSS WL0[81] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4325 VSS WL0[81] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4326 VSS WL0[81] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4327 VSS WL0[81] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4328 VSS WL0[81] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4329 VSS WL0[81] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4330 VSS WL0[81] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4331 VSS WL0[81] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4332 VSS WL0[81] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4333 VSS WL0[81] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4334 VSS WL0[81] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4335 VSS WL0[81] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4336 VSS WL0[81] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4337 VSS WL0[81] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4338 VSS WL0[81] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4339 VSS WL0[81] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4340 VSS WL0[81] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4341 VSS WL0[81] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4342 VSS WL0[81] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4343 VSS WL0[81] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4344 VSS WL0[81] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4345 VSS WL0[81] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4346 VSS WL0[81] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4347 VSS WL0[81] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4348 VSS WL0[81] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4349 VSS WL0[81] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4350 VSS WL0[81] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4351 VSS WL0[81] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4352 VSS WL0[81] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x520
XM4353 VSS WL0[82] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4354 VSS WL0[82] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4355 VSS WL0[82] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4356 VSS WL0[82] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4357 VSS WL0[82] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4358 VSS WL0[82] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4359 VSS WL0[82] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4360 VSS WL0[82] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4361 VSS WL0[82] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4362 VSS WL0[82] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4363 VSS WL0[82] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4364 VSS WL0[82] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4365 VSS WL0[82] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4366 VSS WL0[82] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4367 VSS WL0[82] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4368 VSS WL0[82] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4369 VSS WL0[82] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4370 VSS WL0[82] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4371 VSS WL0[82] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4372 VSS WL0[82] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4373 VSS WL0[82] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4374 VSS WL0[82] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4375 VSS WL0[82] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4376 VSS WL0[82] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4377 VSS WL0[82] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4378 VSS WL0[82] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4379 VSS WL0[82] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4380 VSS WL0[82] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4381 VSS WL0[82] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4382 VSS WL0[82] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4383 VSS WL0[82] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4384 VSS WL0[82] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4385 VSS WL0[82] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4386 VSS WL0[82] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4387 VSS WL0[82] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4388 VSS WL0[82] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4389 VSS WL0[82] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4390 VSS WL0[82] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4391 VSS WL0[82] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4392 VSS WL0[82] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4393 VSS WL0[82] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4394 VSS WL0[82] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4395 VSS WL0[82] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4396 VSS WL0[82] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4397 VSS WL0[82] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4398 VSS WL0[82] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4399 VSS WL0[82] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4400 VSS WL0[82] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4401 VSS WL0[82] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4402 VSS WL0[82] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4403 VSS WL0[82] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4404 VSS WL0[82] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4405 VSS WL0[82] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4406 VSS WL0[82] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4407 VSS WL0[82] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x530
XM4408 VSS WL0[83] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4409 VSS WL0[83] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4410 VSS WL0[83] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4411 VSS WL0[83] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4412 VSS WL0[83] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4413 VSS WL0[83] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4414 VSS WL0[83] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4415 VSS WL0[83] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4416 VSS WL0[83] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4417 VSS WL0[83] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4418 VSS WL0[83] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4419 VSS WL0[83] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4420 VSS WL0[83] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4421 VSS WL0[83] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4422 VSS WL0[83] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4423 VSS WL0[83] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4424 VSS WL0[83] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4425 VSS WL0[83] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4426 VSS WL0[83] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4427 VSS WL0[83] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4428 VSS WL0[83] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4429 VSS WL0[83] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4430 VSS WL0[83] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4431 VSS WL0[83] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4432 VSS WL0[83] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4433 VSS WL0[83] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4434 VSS WL0[83] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4435 VSS WL0[83] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4436 VSS WL0[83] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4437 VSS WL0[83] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4438 VSS WL0[83] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4439 VSS WL0[83] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4440 VSS WL0[83] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4441 VSS WL0[83] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4442 VSS WL0[83] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4443 VSS WL0[83] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4444 VSS WL0[83] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4445 VSS WL0[83] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4446 VSS WL0[83] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4447 VSS WL0[83] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4448 VSS WL0[83] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4449 VSS WL0[83] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4450 VSS WL0[83] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4451 VSS WL0[83] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4452 VSS WL0[83] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4453 VSS WL0[83] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4454 VSS WL0[83] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4455 VSS WL0[83] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4456 VSS WL0[83] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4457 VSS WL0[83] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4458 VSS WL0[83] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4459 VSS WL0[83] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4460 VSS WL0[83] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4461 VSS WL0[83] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x540
XM4462 VSS WL0[84] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4463 VSS WL0[84] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4464 VSS WL0[84] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4465 VSS WL0[84] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4466 VSS WL0[84] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4467 VSS WL0[84] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4468 VSS WL0[84] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4469 VSS WL0[84] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4470 VSS WL0[84] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4471 VSS WL0[84] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4472 VSS WL0[84] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4473 VSS WL0[84] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4474 VSS WL0[84] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4475 VSS WL0[84] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4476 VSS WL0[84] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4477 VSS WL0[84] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4478 VSS WL0[84] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4479 VSS WL0[84] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4480 VSS WL0[84] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4481 VSS WL0[84] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4482 VSS WL0[84] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4483 VSS WL0[84] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4484 VSS WL0[84] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4485 VSS WL0[84] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4486 VSS WL0[84] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4487 VSS WL0[84] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4488 VSS WL0[84] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4489 VSS WL0[84] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4490 VSS WL0[84] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4491 VSS WL0[84] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4492 VSS WL0[84] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4493 VSS WL0[84] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4494 VSS WL0[84] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4495 VSS WL0[84] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4496 VSS WL0[84] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4497 VSS WL0[84] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4498 VSS WL0[84] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4499 VSS WL0[84] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4500 VSS WL0[84] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4501 VSS WL0[84] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4502 VSS WL0[84] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4503 VSS WL0[84] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4504 VSS WL0[84] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4505 VSS WL0[84] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4506 VSS WL0[84] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4507 VSS WL0[84] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4508 VSS WL0[84] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4509 VSS WL0[84] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4510 VSS WL0[84] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4511 VSS WL0[84] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4512 VSS WL0[84] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4513 VSS WL0[84] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4514 VSS WL0[84] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4515 VSS WL0[84] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4516 VSS WL0[84] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4517 VSS WL0[84] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4518 VSS WL0[84] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4519 VSS WL0[84] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4520 VSS WL0[84] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4521 VSS WL0[84] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4522 VSS WL0[84] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4523 VSS WL0[84] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x550
XM4524 VSS WL0[85] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4525 VSS WL0[85] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4526 VSS WL0[85] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4527 VSS WL0[85] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4528 VSS WL0[85] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4529 VSS WL0[85] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4530 VSS WL0[85] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4531 VSS WL0[85] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4532 VSS WL0[85] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4533 VSS WL0[85] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4534 VSS WL0[85] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4535 VSS WL0[85] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4536 VSS WL0[85] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4537 VSS WL0[85] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4538 VSS WL0[85] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4539 VSS WL0[85] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4540 VSS WL0[85] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4541 VSS WL0[85] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4542 VSS WL0[85] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4543 VSS WL0[85] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4544 VSS WL0[85] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4545 VSS WL0[85] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4546 VSS WL0[85] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4547 VSS WL0[85] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4548 VSS WL0[85] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4549 VSS WL0[85] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4550 VSS WL0[85] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4551 VSS WL0[85] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4552 VSS WL0[85] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4553 VSS WL0[85] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4554 VSS WL0[85] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4555 VSS WL0[85] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4556 VSS WL0[85] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4557 VSS WL0[85] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4558 VSS WL0[85] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4559 VSS WL0[85] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4560 VSS WL0[85] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4561 VSS WL0[85] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4562 VSS WL0[85] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4563 VSS WL0[85] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4564 VSS WL0[85] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4565 VSS WL0[85] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4566 VSS WL0[85] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4567 VSS WL0[85] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4568 VSS WL0[85] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4569 VSS WL0[85] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4570 VSS WL0[85] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4571 VSS WL0[85] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4572 VSS WL0[85] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4573 VSS WL0[85] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x560
XM4574 VSS WL0[86] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4575 VSS WL0[86] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4576 VSS WL0[86] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4577 VSS WL0[86] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4578 VSS WL0[86] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4579 VSS WL0[86] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4580 VSS WL0[86] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4581 VSS WL0[86] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4582 VSS WL0[86] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4583 VSS WL0[86] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4584 VSS WL0[86] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4585 VSS WL0[86] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4586 VSS WL0[86] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4587 VSS WL0[86] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4588 VSS WL0[86] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4589 VSS WL0[86] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4590 VSS WL0[86] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4591 VSS WL0[86] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4592 VSS WL0[86] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4593 VSS WL0[86] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4594 VSS WL0[86] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4595 VSS WL0[86] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4596 VSS WL0[86] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4597 VSS WL0[86] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4598 VSS WL0[86] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4599 VSS WL0[86] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4600 VSS WL0[86] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4601 VSS WL0[86] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4602 VSS WL0[86] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4603 VSS WL0[86] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4604 VSS WL0[86] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4605 VSS WL0[86] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4606 VSS WL0[86] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4607 VSS WL0[86] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4608 VSS WL0[86] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4609 VSS WL0[86] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4610 VSS WL0[86] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4611 VSS WL0[86] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4612 VSS WL0[86] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4613 VSS WL0[86] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4614 VSS WL0[86] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4615 VSS WL0[86] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4616 VSS WL0[86] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4617 VSS WL0[86] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4618 VSS WL0[86] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4619 VSS WL0[86] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4620 VSS WL0[86] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4621 VSS WL0[86] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4622 VSS WL0[86] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4623 VSS WL0[86] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4624 VSS WL0[86] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4625 VSS WL0[86] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4626 VSS WL0[86] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4627 VSS WL0[86] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4628 VSS WL0[86] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4629 VSS WL0[86] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4630 VSS WL0[86] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4631 VSS WL0[86] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4632 VSS WL0[86] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4633 VSS WL0[86] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4634 VSS WL0[86] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4635 VSS WL0[86] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4636 VSS WL0[86] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4637 VSS WL0[86] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4638 VSS WL0[86] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4639 VSS WL0[86] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4640 VSS WL0[86] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4641 VSS WL0[86] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4642 VSS WL0[86] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4643 VSS WL0[86] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4644 VSS WL0[86] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4645 VSS WL0[86] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4646 VSS WL0[86] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x570
XM4647 VSS WL0[87] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4648 VSS WL0[87] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4649 VSS WL0[87] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4650 VSS WL0[87] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4651 VSS WL0[87] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4652 VSS WL0[87] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4653 VSS WL0[87] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4654 VSS WL0[87] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4655 VSS WL0[87] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4656 VSS WL0[87] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4657 VSS WL0[87] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4658 VSS WL0[87] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4659 VSS WL0[87] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4660 VSS WL0[87] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4661 VSS WL0[87] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4662 VSS WL0[87] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4663 VSS WL0[87] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4664 VSS WL0[87] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4665 VSS WL0[87] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4666 VSS WL0[87] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4667 VSS WL0[87] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4668 VSS WL0[87] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4669 VSS WL0[87] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4670 VSS WL0[87] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4671 VSS WL0[87] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4672 VSS WL0[87] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4673 VSS WL0[87] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4674 VSS WL0[87] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4675 VSS WL0[87] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4676 VSS WL0[87] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4677 VSS WL0[87] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4678 VSS WL0[87] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4679 VSS WL0[87] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4680 VSS WL0[87] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4681 VSS WL0[87] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4682 VSS WL0[87] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4683 VSS WL0[87] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4684 VSS WL0[87] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4685 VSS WL0[87] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4686 VSS WL0[87] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4687 VSS WL0[87] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4688 VSS WL0[87] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4689 VSS WL0[87] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4690 VSS WL0[87] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4691 VSS WL0[87] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4692 VSS WL0[87] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4693 VSS WL0[87] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4694 VSS WL0[87] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4695 VSS WL0[87] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4696 VSS WL0[87] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x580
XM4697 VSS WL0[88] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4698 VSS WL0[88] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4699 VSS WL0[88] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4700 VSS WL0[88] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4701 VSS WL0[88] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4702 VSS WL0[88] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4703 VSS WL0[88] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4704 VSS WL0[88] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4705 VSS WL0[88] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4706 VSS WL0[88] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4707 VSS WL0[88] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4708 VSS WL0[88] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4709 VSS WL0[88] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4710 VSS WL0[88] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4711 VSS WL0[88] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4712 VSS WL0[88] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4713 VSS WL0[88] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4714 VSS WL0[88] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4715 VSS WL0[88] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4716 VSS WL0[88] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4717 VSS WL0[88] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4718 VSS WL0[88] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4719 VSS WL0[88] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4720 VSS WL0[88] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4721 VSS WL0[88] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4722 VSS WL0[88] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4723 VSS WL0[88] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4724 VSS WL0[88] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4725 VSS WL0[88] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4726 VSS WL0[88] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4727 VSS WL0[88] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4728 VSS WL0[88] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4729 VSS WL0[88] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4730 VSS WL0[88] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4731 VSS WL0[88] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4732 VSS WL0[88] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4733 VSS WL0[88] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4734 VSS WL0[88] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4735 VSS WL0[88] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4736 VSS WL0[88] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4737 VSS WL0[88] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x590
XM4738 VSS WL0[89] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4739 VSS WL0[89] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4740 VSS WL0[89] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4741 VSS WL0[89] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4742 VSS WL0[89] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4743 VSS WL0[89] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4744 VSS WL0[89] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4745 VSS WL0[89] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4746 VSS WL0[89] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4747 VSS WL0[89] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4748 VSS WL0[89] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4749 VSS WL0[89] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4750 VSS WL0[89] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4751 VSS WL0[89] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4752 VSS WL0[89] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4753 VSS WL0[89] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4754 VSS WL0[89] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4755 VSS WL0[89] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4756 VSS WL0[89] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4757 VSS WL0[89] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4758 VSS WL0[89] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4759 VSS WL0[89] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4760 VSS WL0[89] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4761 VSS WL0[89] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4762 VSS WL0[89] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4763 VSS WL0[89] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4764 VSS WL0[89] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4765 VSS WL0[89] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4766 VSS WL0[89] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4767 VSS WL0[89] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4768 VSS WL0[89] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4769 VSS WL0[89] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4770 VSS WL0[89] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4771 VSS WL0[89] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4772 VSS WL0[89] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4773 VSS WL0[89] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4774 VSS WL0[89] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4775 VSS WL0[89] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4776 VSS WL0[89] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4777 VSS WL0[89] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4778 VSS WL0[89] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4779 VSS WL0[89] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4780 VSS WL0[89] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4781 VSS WL0[89] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4782 VSS WL0[89] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4783 VSS WL0[89] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4784 VSS WL0[89] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4785 VSS WL0[89] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4786 VSS WL0[89] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4787 VSS WL0[89] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x5a0
XM4788 VSS WL0[90] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4789 VSS WL0[90] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4790 VSS WL0[90] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4791 VSS WL0[90] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4792 VSS WL0[90] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4793 VSS WL0[90] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4794 VSS WL0[90] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4795 VSS WL0[90] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4796 VSS WL0[90] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4797 VSS WL0[90] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4798 VSS WL0[90] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4799 VSS WL0[90] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4800 VSS WL0[90] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4801 VSS WL0[90] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4802 VSS WL0[90] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4803 VSS WL0[90] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4804 VSS WL0[90] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4805 VSS WL0[90] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4806 VSS WL0[90] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4807 VSS WL0[90] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4808 VSS WL0[90] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4809 VSS WL0[90] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4810 VSS WL0[90] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4811 VSS WL0[90] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4812 VSS WL0[90] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4813 VSS WL0[90] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4814 VSS WL0[90] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4815 VSS WL0[90] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4816 VSS WL0[90] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4817 VSS WL0[90] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4818 VSS WL0[90] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4819 VSS WL0[90] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4820 VSS WL0[90] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4821 VSS WL0[90] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4822 VSS WL0[90] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4823 VSS WL0[90] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4824 VSS WL0[90] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4825 VSS WL0[90] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4826 VSS WL0[90] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4827 VSS WL0[90] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4828 VSS WL0[90] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4829 VSS WL0[90] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4830 VSS WL0[90] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4831 VSS WL0[90] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4832 VSS WL0[90] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4833 VSS WL0[90] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4834 VSS WL0[90] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4835 VSS WL0[90] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4836 VSS WL0[90] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4837 VSS WL0[90] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4838 VSS WL0[90] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4839 VSS WL0[90] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4840 VSS WL0[90] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4841 VSS WL0[90] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x5b0
XM4842 VSS WL0[91] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4843 VSS WL0[91] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4844 VSS WL0[91] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4845 VSS WL0[91] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4846 VSS WL0[91] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4847 VSS WL0[91] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4848 VSS WL0[91] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4849 VSS WL0[91] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4850 VSS WL0[91] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4851 VSS WL0[91] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4852 VSS WL0[91] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4853 VSS WL0[91] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4854 VSS WL0[91] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4855 VSS WL0[91] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4856 VSS WL0[91] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4857 VSS WL0[91] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4858 VSS WL0[91] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4859 VSS WL0[91] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4860 VSS WL0[91] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4861 VSS WL0[91] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4862 VSS WL0[91] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4863 VSS WL0[91] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4864 VSS WL0[91] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4865 VSS WL0[91] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4866 VSS WL0[91] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4867 VSS WL0[91] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4868 VSS WL0[91] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4869 VSS WL0[91] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4870 VSS WL0[91] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4871 VSS WL0[91] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4872 VSS WL0[91] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4873 VSS WL0[91] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4874 VSS WL0[91] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4875 VSS WL0[91] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4876 VSS WL0[91] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4877 VSS WL0[91] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x5c0
XM4878 VSS WL0[92] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4879 VSS WL0[92] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4880 VSS WL0[92] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4881 VSS WL0[92] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4882 VSS WL0[92] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4883 VSS WL0[92] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4884 VSS WL0[92] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4885 VSS WL0[92] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4886 VSS WL0[92] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4887 VSS WL0[92] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4888 VSS WL0[92] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4889 VSS WL0[92] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4890 VSS WL0[92] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4891 VSS WL0[92] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4892 VSS WL0[92] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4893 VSS WL0[92] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4894 VSS WL0[92] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4895 VSS WL0[92] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4896 VSS WL0[92] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4897 VSS WL0[92] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4898 VSS WL0[92] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4899 VSS WL0[92] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4900 VSS WL0[92] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4901 VSS WL0[92] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4902 VSS WL0[92] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4903 VSS WL0[92] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4904 VSS WL0[92] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4905 VSS WL0[92] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4906 VSS WL0[92] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4907 VSS WL0[92] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4908 VSS WL0[92] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4909 VSS WL0[92] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4910 VSS WL0[92] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4911 VSS WL0[92] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4912 VSS WL0[92] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4913 VSS WL0[92] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4914 VSS WL0[92] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4915 VSS WL0[92] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4916 VSS WL0[92] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4917 VSS WL0[92] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4918 VSS WL0[92] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4919 VSS WL0[92] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4920 VSS WL0[92] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4921 VSS WL0[92] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4922 VSS WL0[92] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4923 VSS WL0[92] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4924 VSS WL0[92] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4925 VSS WL0[92] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4926 VSS WL0[92] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4927 VSS WL0[92] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4928 VSS WL0[92] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4929 VSS WL0[92] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4930 VSS WL0[92] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x5d0
XM4931 VSS WL0[93] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4932 VSS WL0[93] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4933 VSS WL0[93] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4934 VSS WL0[93] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4935 VSS WL0[93] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4936 VSS WL0[93] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4937 VSS WL0[93] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4938 VSS WL0[93] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4939 VSS WL0[93] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4940 VSS WL0[93] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4941 VSS WL0[93] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4942 VSS WL0[93] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4943 VSS WL0[93] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4944 VSS WL0[93] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4945 VSS WL0[93] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4946 VSS WL0[93] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4947 VSS WL0[93] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4948 VSS WL0[93] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4949 VSS WL0[93] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4950 VSS WL0[93] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4951 VSS WL0[93] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4952 VSS WL0[93] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4953 VSS WL0[93] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4954 VSS WL0[93] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4955 VSS WL0[93] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4956 VSS WL0[93] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4957 VSS WL0[93] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4958 VSS WL0[93] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4959 VSS WL0[93] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4960 VSS WL0[93] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4961 VSS WL0[93] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4962 VSS WL0[93] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4963 VSS WL0[93] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4964 VSS WL0[93] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4965 VSS WL0[93] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4966 VSS WL0[93] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4967 VSS WL0[93] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4968 VSS WL0[93] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4969 VSS WL0[93] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4970 VSS WL0[93] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4971 VSS WL0[93] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4972 VSS WL0[93] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4973 VSS WL0[93] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4974 VSS WL0[93] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x5e0
XM4975 VSS WL0[94] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4976 VSS WL0[94] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4977 VSS WL0[94] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4978 VSS WL0[94] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4979 VSS WL0[94] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4980 VSS WL0[94] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4981 VSS WL0[94] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4982 VSS WL0[94] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4983 VSS WL0[94] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4984 VSS WL0[94] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4985 VSS WL0[94] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4986 VSS WL0[94] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4987 VSS WL0[94] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4988 VSS WL0[94] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4989 VSS WL0[94] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4990 VSS WL0[94] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4991 VSS WL0[94] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4992 VSS WL0[94] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4993 VSS WL0[94] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4994 VSS WL0[94] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4995 VSS WL0[94] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4996 VSS WL0[94] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4997 VSS WL0[94] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4998 VSS WL0[94] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM4999 VSS WL0[94] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5000 VSS WL0[94] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5001 VSS WL0[94] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5002 VSS WL0[94] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5003 VSS WL0[94] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5004 VSS WL0[94] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5005 VSS WL0[94] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5006 VSS WL0[94] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5007 VSS WL0[94] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5008 VSS WL0[94] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5009 VSS WL0[94] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5010 VSS WL0[94] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5011 VSS WL0[94] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5012 VSS WL0[94] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5013 VSS WL0[94] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5014 VSS WL0[94] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5015 VSS WL0[94] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5016 VSS WL0[94] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5017 VSS WL0[94] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5018 VSS WL0[94] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5019 VSS WL0[94] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5020 VSS WL0[94] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5021 VSS WL0[94] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5022 VSS WL0[94] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5023 VSS WL0[94] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5024 VSS WL0[94] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5025 VSS WL0[94] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5026 VSS WL0[94] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x5f0
XM5027 VSS WL0[95] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5028 VSS WL0[95] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5029 VSS WL0[95] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5030 VSS WL0[95] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5031 VSS WL0[95] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5032 VSS WL0[95] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5033 VSS WL0[95] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5034 VSS WL0[95] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5035 VSS WL0[95] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5036 VSS WL0[95] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5037 VSS WL0[95] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5038 VSS WL0[95] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5039 VSS WL0[95] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5040 VSS WL0[95] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5041 VSS WL0[95] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5042 VSS WL0[95] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5043 VSS WL0[95] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5044 VSS WL0[95] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5045 VSS WL0[95] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5046 VSS WL0[95] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5047 VSS WL0[95] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5048 VSS WL0[95] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5049 VSS WL0[95] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5050 VSS WL0[95] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5051 VSS WL0[95] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5052 VSS WL0[95] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5053 VSS WL0[95] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5054 VSS WL0[95] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5055 VSS WL0[95] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5056 VSS WL0[95] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5057 VSS WL0[95] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5058 VSS WL0[95] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5059 VSS WL0[95] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5060 VSS WL0[95] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5061 VSS WL0[95] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5062 VSS WL0[95] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5063 VSS WL0[95] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5064 VSS WL0[95] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5065 VSS WL0[95] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5066 VSS WL0[95] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5067 VSS WL0[95] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5068 VSS WL0[95] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5069 VSS WL0[95] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5070 VSS WL0[95] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5071 VSS WL0[95] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x600
XM5072 VSS WL0[96] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5073 VSS WL0[96] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5074 VSS WL0[96] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5075 VSS WL0[96] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5076 VSS WL0[96] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5077 VSS WL0[96] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5078 VSS WL0[96] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5079 VSS WL0[96] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5080 VSS WL0[96] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5081 VSS WL0[96] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5082 VSS WL0[96] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5083 VSS WL0[96] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5084 VSS WL0[96] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5085 VSS WL0[96] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5086 VSS WL0[96] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5087 VSS WL0[96] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5088 VSS WL0[96] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5089 VSS WL0[96] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5090 VSS WL0[96] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5091 VSS WL0[96] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5092 VSS WL0[96] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5093 VSS WL0[96] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5094 VSS WL0[96] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5095 VSS WL0[96] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5096 VSS WL0[96] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5097 VSS WL0[96] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5098 VSS WL0[96] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5099 VSS WL0[96] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5100 VSS WL0[96] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5101 VSS WL0[96] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5102 VSS WL0[96] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5103 VSS WL0[96] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5104 VSS WL0[96] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5105 VSS WL0[96] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5106 VSS WL0[96] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5107 VSS WL0[96] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5108 VSS WL0[96] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5109 VSS WL0[96] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5110 VSS WL0[96] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5111 VSS WL0[96] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5112 VSS WL0[96] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5113 VSS WL0[96] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5114 VSS WL0[96] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5115 VSS WL0[96] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x610
XM5116 VSS WL0[97] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5117 VSS WL0[97] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5118 VSS WL0[97] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5119 VSS WL0[97] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5120 VSS WL0[97] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5121 VSS WL0[97] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5122 VSS WL0[97] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5123 VSS WL0[97] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5124 VSS WL0[97] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5125 VSS WL0[97] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5126 VSS WL0[97] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5127 VSS WL0[97] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5128 VSS WL0[97] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5129 VSS WL0[97] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5130 VSS WL0[97] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5131 VSS WL0[97] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5132 VSS WL0[97] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5133 VSS WL0[97] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5134 VSS WL0[97] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5135 VSS WL0[97] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5136 VSS WL0[97] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5137 VSS WL0[97] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5138 VSS WL0[97] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5139 VSS WL0[97] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5140 VSS WL0[97] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5141 VSS WL0[97] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5142 VSS WL0[97] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5143 VSS WL0[97] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5144 VSS WL0[97] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5145 VSS WL0[97] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5146 VSS WL0[97] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5147 VSS WL0[97] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5148 VSS WL0[97] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5149 VSS WL0[97] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5150 VSS WL0[97] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5151 VSS WL0[97] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5152 VSS WL0[97] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5153 VSS WL0[97] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5154 VSS WL0[97] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5155 VSS WL0[97] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5156 VSS WL0[97] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5157 VSS WL0[97] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5158 VSS WL0[97] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5159 VSS WL0[97] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5160 VSS WL0[97] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5161 VSS WL0[97] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5162 VSS WL0[97] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5163 VSS WL0[97] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5164 VSS WL0[97] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5165 VSS WL0[97] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5166 VSS WL0[97] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5167 VSS WL0[97] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5168 VSS WL0[97] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x620
XM5169 VSS WL0[98] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5170 VSS WL0[98] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5171 VSS WL0[98] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5172 VSS WL0[98] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5173 VSS WL0[98] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5174 VSS WL0[98] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5175 VSS WL0[98] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5176 VSS WL0[98] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5177 VSS WL0[98] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5178 VSS WL0[98] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5179 VSS WL0[98] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5180 VSS WL0[98] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5181 VSS WL0[98] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5182 VSS WL0[98] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5183 VSS WL0[98] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5184 VSS WL0[98] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5185 VSS WL0[98] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5186 VSS WL0[98] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5187 VSS WL0[98] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5188 VSS WL0[98] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5189 VSS WL0[98] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5190 VSS WL0[98] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5191 VSS WL0[98] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5192 VSS WL0[98] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5193 VSS WL0[98] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5194 VSS WL0[98] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5195 VSS WL0[98] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5196 VSS WL0[98] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5197 VSS WL0[98] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5198 VSS WL0[98] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5199 VSS WL0[98] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5200 VSS WL0[98] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5201 VSS WL0[98] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5202 VSS WL0[98] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5203 VSS WL0[98] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5204 VSS WL0[98] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5205 VSS WL0[98] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5206 VSS WL0[98] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5207 VSS WL0[98] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5208 VSS WL0[98] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5209 VSS WL0[98] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5210 VSS WL0[98] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x630
XM5211 VSS WL0[99] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5212 VSS WL0[99] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5213 VSS WL0[99] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5214 VSS WL0[99] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5215 VSS WL0[99] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5216 VSS WL0[99] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5217 VSS WL0[99] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5218 VSS WL0[99] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5219 VSS WL0[99] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5220 VSS WL0[99] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5221 VSS WL0[99] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5222 VSS WL0[99] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5223 VSS WL0[99] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5224 VSS WL0[99] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5225 VSS WL0[99] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5226 VSS WL0[99] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5227 VSS WL0[99] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5228 VSS WL0[99] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5229 VSS WL0[99] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5230 VSS WL0[99] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5231 VSS WL0[99] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5232 VSS WL0[99] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5233 VSS WL0[99] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5234 VSS WL0[99] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5235 VSS WL0[99] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5236 VSS WL0[99] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5237 VSS WL0[99] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5238 VSS WL0[99] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5239 VSS WL0[99] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5240 VSS WL0[99] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5241 VSS WL0[99] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5242 VSS WL0[99] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5243 VSS WL0[99] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5244 VSS WL0[99] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5245 VSS WL0[99] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5246 VSS WL0[99] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5247 VSS WL0[99] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5248 VSS WL0[99] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5249 VSS WL0[99] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5250 VSS WL0[99] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5251 VSS WL0[99] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5252 VSS WL0[99] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5253 VSS WL0[99] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5254 VSS WL0[99] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5255 VSS WL0[99] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5256 VSS WL0[99] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5257 VSS WL0[99] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5258 VSS WL0[99] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5259 VSS WL0[99] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5260 VSS WL0[99] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5261 VSS WL0[99] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5262 VSS WL0[99] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5263 VSS WL0[99] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5264 VSS WL0[99] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5265 VSS WL0[99] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5266 VSS WL0[99] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5267 VSS WL0[99] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5268 VSS WL0[99] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5269 VSS WL0[99] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5270 VSS WL0[99] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5271 VSS WL0[99] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5272 VSS WL0[99] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5273 VSS WL0[99] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x640
XM5274 VSS WL0[100] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5275 VSS WL0[100] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5276 VSS WL0[100] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5277 VSS WL0[100] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5278 VSS WL0[100] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5279 VSS WL0[100] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5280 VSS WL0[100] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5281 VSS WL0[100] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5282 VSS WL0[100] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5283 VSS WL0[100] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5284 VSS WL0[100] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5285 VSS WL0[100] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5286 VSS WL0[100] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5287 VSS WL0[100] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5288 VSS WL0[100] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5289 VSS WL0[100] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5290 VSS WL0[100] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5291 VSS WL0[100] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5292 VSS WL0[100] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5293 VSS WL0[100] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5294 VSS WL0[100] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5295 VSS WL0[100] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5296 VSS WL0[100] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5297 VSS WL0[100] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5298 VSS WL0[100] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5299 VSS WL0[100] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5300 VSS WL0[100] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5301 VSS WL0[100] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5302 VSS WL0[100] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5303 VSS WL0[100] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5304 VSS WL0[100] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5305 VSS WL0[100] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5306 VSS WL0[100] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5307 VSS WL0[100] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5308 VSS WL0[100] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5309 VSS WL0[100] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5310 VSS WL0[100] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5311 VSS WL0[100] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5312 VSS WL0[100] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5313 VSS WL0[100] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5314 VSS WL0[100] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5315 VSS WL0[100] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5316 VSS WL0[100] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5317 VSS WL0[100] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5318 VSS WL0[100] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5319 VSS WL0[100] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5320 VSS WL0[100] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5321 VSS WL0[100] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5322 VSS WL0[100] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5323 VSS WL0[100] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5324 VSS WL0[100] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5325 VSS WL0[100] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5326 VSS WL0[100] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x650
XM5327 VSS WL0[101] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5328 VSS WL0[101] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5329 VSS WL0[101] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5330 VSS WL0[101] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5331 VSS WL0[101] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5332 VSS WL0[101] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5333 VSS WL0[101] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5334 VSS WL0[101] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5335 VSS WL0[101] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5336 VSS WL0[101] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5337 VSS WL0[101] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5338 VSS WL0[101] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5339 VSS WL0[101] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5340 VSS WL0[101] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5341 VSS WL0[101] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5342 VSS WL0[101] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5343 VSS WL0[101] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5344 VSS WL0[101] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5345 VSS WL0[101] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5346 VSS WL0[101] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5347 VSS WL0[101] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5348 VSS WL0[101] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5349 VSS WL0[101] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5350 VSS WL0[101] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5351 VSS WL0[101] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5352 VSS WL0[101] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5353 VSS WL0[101] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5354 VSS WL0[101] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5355 VSS WL0[101] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5356 VSS WL0[101] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5357 VSS WL0[101] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5358 VSS WL0[101] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5359 VSS WL0[101] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5360 VSS WL0[101] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5361 VSS WL0[101] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5362 VSS WL0[101] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5363 VSS WL0[101] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5364 VSS WL0[101] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5365 VSS WL0[101] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5366 VSS WL0[101] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5367 VSS WL0[101] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5368 VSS WL0[101] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5369 VSS WL0[101] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5370 VSS WL0[101] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5371 VSS WL0[101] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5372 VSS WL0[101] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5373 VSS WL0[101] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5374 VSS WL0[101] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5375 VSS WL0[101] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5376 VSS WL0[101] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5377 VSS WL0[101] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5378 VSS WL0[101] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5379 VSS WL0[101] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5380 VSS WL0[101] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5381 VSS WL0[101] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5382 VSS WL0[101] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5383 VSS WL0[101] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5384 VSS WL0[101] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5385 VSS WL0[101] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5386 VSS WL0[101] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5387 VSS WL0[101] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5388 VSS WL0[101] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5389 VSS WL0[101] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5390 VSS WL0[101] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5391 VSS WL0[101] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5392 VSS WL0[101] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5393 VSS WL0[101] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5394 VSS WL0[101] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5395 VSS WL0[101] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5396 VSS WL0[101] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5397 VSS WL0[101] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5398 VSS WL0[101] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5399 VSS WL0[101] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5400 VSS WL0[101] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5401 VSS WL0[101] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5402 VSS WL0[101] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x660
XM5403 VSS WL0[102] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5404 VSS WL0[102] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5405 VSS WL0[102] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5406 VSS WL0[102] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5407 VSS WL0[102] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5408 VSS WL0[102] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5409 VSS WL0[102] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5410 VSS WL0[102] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5411 VSS WL0[102] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5412 VSS WL0[102] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5413 VSS WL0[102] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5414 VSS WL0[102] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5415 VSS WL0[102] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5416 VSS WL0[102] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5417 VSS WL0[102] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5418 VSS WL0[102] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5419 VSS WL0[102] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5420 VSS WL0[102] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5421 VSS WL0[102] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5422 VSS WL0[102] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5423 VSS WL0[102] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5424 VSS WL0[102] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5425 VSS WL0[102] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5426 VSS WL0[102] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5427 VSS WL0[102] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5428 VSS WL0[102] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5429 VSS WL0[102] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5430 VSS WL0[102] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5431 VSS WL0[102] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5432 VSS WL0[102] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5433 VSS WL0[102] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5434 VSS WL0[102] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5435 VSS WL0[102] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5436 VSS WL0[102] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5437 VSS WL0[102] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5438 VSS WL0[102] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5439 VSS WL0[102] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5440 VSS WL0[102] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5441 VSS WL0[102] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5442 VSS WL0[102] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5443 VSS WL0[102] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5444 VSS WL0[102] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5445 VSS WL0[102] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5446 VSS WL0[102] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5447 VSS WL0[102] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5448 VSS WL0[102] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5449 VSS WL0[102] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5450 VSS WL0[102] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5451 VSS WL0[102] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5452 VSS WL0[102] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5453 VSS WL0[102] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5454 VSS WL0[102] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5455 VSS WL0[102] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5456 VSS WL0[102] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5457 VSS WL0[102] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5458 VSS WL0[102] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5459 VSS WL0[102] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5460 VSS WL0[102] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x670
XM5461 VSS WL0[103] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5462 VSS WL0[103] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5463 VSS WL0[103] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5464 VSS WL0[103] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5465 VSS WL0[103] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5466 VSS WL0[103] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5467 VSS WL0[103] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5468 VSS WL0[103] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5469 VSS WL0[103] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5470 VSS WL0[103] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5471 VSS WL0[103] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5472 VSS WL0[103] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5473 VSS WL0[103] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5474 VSS WL0[103] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5475 VSS WL0[103] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5476 VSS WL0[103] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5477 VSS WL0[103] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5478 VSS WL0[103] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5479 VSS WL0[103] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5480 VSS WL0[103] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5481 VSS WL0[103] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5482 VSS WL0[103] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5483 VSS WL0[103] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5484 VSS WL0[103] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5485 VSS WL0[103] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5486 VSS WL0[103] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5487 VSS WL0[103] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5488 VSS WL0[103] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5489 VSS WL0[103] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5490 VSS WL0[103] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5491 VSS WL0[103] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5492 VSS WL0[103] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5493 VSS WL0[103] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5494 VSS WL0[103] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5495 VSS WL0[103] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5496 VSS WL0[103] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5497 VSS WL0[103] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5498 VSS WL0[103] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5499 VSS WL0[103] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5500 VSS WL0[103] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5501 VSS WL0[103] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5502 VSS WL0[103] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5503 VSS WL0[103] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5504 VSS WL0[103] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5505 VSS WL0[103] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5506 VSS WL0[103] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x680
XM5507 VSS WL0[104] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5508 VSS WL0[104] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5509 VSS WL0[104] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5510 VSS WL0[104] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5511 VSS WL0[104] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5512 VSS WL0[104] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5513 VSS WL0[104] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5514 VSS WL0[104] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5515 VSS WL0[104] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5516 VSS WL0[104] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5517 VSS WL0[104] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5518 VSS WL0[104] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5519 VSS WL0[104] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5520 VSS WL0[104] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5521 VSS WL0[104] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5522 VSS WL0[104] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5523 VSS WL0[104] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5524 VSS WL0[104] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5525 VSS WL0[104] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5526 VSS WL0[104] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5527 VSS WL0[104] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5528 VSS WL0[104] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5529 VSS WL0[104] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5530 VSS WL0[104] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5531 VSS WL0[104] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5532 VSS WL0[104] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5533 VSS WL0[104] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5534 VSS WL0[104] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5535 VSS WL0[104] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5536 VSS WL0[104] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5537 VSS WL0[104] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5538 VSS WL0[104] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5539 VSS WL0[104] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5540 VSS WL0[104] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5541 VSS WL0[104] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5542 VSS WL0[104] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5543 VSS WL0[104] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5544 VSS WL0[104] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5545 VSS WL0[104] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5546 VSS WL0[104] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5547 VSS WL0[104] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5548 VSS WL0[104] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5549 VSS WL0[104] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5550 VSS WL0[104] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5551 VSS WL0[104] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5552 VSS WL0[104] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5553 VSS WL0[104] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5554 VSS WL0[104] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5555 VSS WL0[104] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5556 VSS WL0[104] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x690
XM5557 VSS WL0[105] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5558 VSS WL0[105] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5559 VSS WL0[105] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5560 VSS WL0[105] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5561 VSS WL0[105] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5562 VSS WL0[105] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5563 VSS WL0[105] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5564 VSS WL0[105] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5565 VSS WL0[105] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5566 VSS WL0[105] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5567 VSS WL0[105] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5568 VSS WL0[105] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5569 VSS WL0[105] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5570 VSS WL0[105] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5571 VSS WL0[105] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5572 VSS WL0[105] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5573 VSS WL0[105] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5574 VSS WL0[105] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5575 VSS WL0[105] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5576 VSS WL0[105] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5577 VSS WL0[105] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5578 VSS WL0[105] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5579 VSS WL0[105] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5580 VSS WL0[105] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5581 VSS WL0[105] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5582 VSS WL0[105] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5583 VSS WL0[105] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5584 VSS WL0[105] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5585 VSS WL0[105] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5586 VSS WL0[105] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5587 VSS WL0[105] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5588 VSS WL0[105] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5589 VSS WL0[105] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5590 VSS WL0[105] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5591 VSS WL0[105] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5592 VSS WL0[105] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5593 VSS WL0[105] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5594 VSS WL0[105] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5595 VSS WL0[105] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5596 VSS WL0[105] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5597 VSS WL0[105] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5598 VSS WL0[105] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5599 VSS WL0[105] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x6a0
XM5600 VSS WL0[106] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5601 VSS WL0[106] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5602 VSS WL0[106] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5603 VSS WL0[106] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5604 VSS WL0[106] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5605 VSS WL0[106] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5606 VSS WL0[106] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5607 VSS WL0[106] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5608 VSS WL0[106] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5609 VSS WL0[106] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5610 VSS WL0[106] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5611 VSS WL0[106] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5612 VSS WL0[106] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5613 VSS WL0[106] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5614 VSS WL0[106] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5615 VSS WL0[106] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5616 VSS WL0[106] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5617 VSS WL0[106] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5618 VSS WL0[106] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5619 VSS WL0[106] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5620 VSS WL0[106] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5621 VSS WL0[106] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5622 VSS WL0[106] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5623 VSS WL0[106] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5624 VSS WL0[106] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5625 VSS WL0[106] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5626 VSS WL0[106] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5627 VSS WL0[106] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5628 VSS WL0[106] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5629 VSS WL0[106] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5630 VSS WL0[106] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5631 VSS WL0[106] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5632 VSS WL0[106] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5633 VSS WL0[106] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5634 VSS WL0[106] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5635 VSS WL0[106] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5636 VSS WL0[106] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5637 VSS WL0[106] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5638 VSS WL0[106] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5639 VSS WL0[106] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5640 VSS WL0[106] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5641 VSS WL0[106] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5642 VSS WL0[106] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5643 VSS WL0[106] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5644 VSS WL0[106] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5645 VSS WL0[106] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5646 VSS WL0[106] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5647 VSS WL0[106] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5648 VSS WL0[106] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5649 VSS WL0[106] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x6b0
XM5650 VSS WL0[107] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5651 VSS WL0[107] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5652 VSS WL0[107] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5653 VSS WL0[107] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5654 VSS WL0[107] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5655 VSS WL0[107] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5656 VSS WL0[107] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5657 VSS WL0[107] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5658 VSS WL0[107] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5659 VSS WL0[107] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5660 VSS WL0[107] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5661 VSS WL0[107] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5662 VSS WL0[107] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5663 VSS WL0[107] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5664 VSS WL0[107] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5665 VSS WL0[107] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5666 VSS WL0[107] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5667 VSS WL0[107] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5668 VSS WL0[107] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5669 VSS WL0[107] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5670 VSS WL0[107] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5671 VSS WL0[107] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5672 VSS WL0[107] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5673 VSS WL0[107] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5674 VSS WL0[107] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5675 VSS WL0[107] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5676 VSS WL0[107] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5677 VSS WL0[107] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5678 VSS WL0[107] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5679 VSS WL0[107] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5680 VSS WL0[107] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5681 VSS WL0[107] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5682 VSS WL0[107] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5683 VSS WL0[107] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5684 VSS WL0[107] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5685 VSS WL0[107] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5686 VSS WL0[107] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5687 VSS WL0[107] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5688 VSS WL0[107] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5689 VSS WL0[107] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5690 VSS WL0[107] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5691 VSS WL0[107] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5692 VSS WL0[107] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5693 VSS WL0[107] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5694 VSS WL0[107] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5695 VSS WL0[107] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5696 VSS WL0[107] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5697 VSS WL0[107] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5698 VSS WL0[107] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5699 VSS WL0[107] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5700 VSS WL0[107] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5701 VSS WL0[107] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5702 VSS WL0[107] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5703 VSS WL0[107] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5704 VSS WL0[107] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5705 VSS WL0[107] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5706 VSS WL0[107] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x6c0
XM5707 VSS WL0[108] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5708 VSS WL0[108] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5709 VSS WL0[108] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5710 VSS WL0[108] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5711 VSS WL0[108] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5712 VSS WL0[108] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5713 VSS WL0[108] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5714 VSS WL0[108] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5715 VSS WL0[108] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5716 VSS WL0[108] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5717 VSS WL0[108] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5718 VSS WL0[108] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5719 VSS WL0[108] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5720 VSS WL0[108] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5721 VSS WL0[108] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5722 VSS WL0[108] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5723 VSS WL0[108] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5724 VSS WL0[108] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5725 VSS WL0[108] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5726 VSS WL0[108] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5727 VSS WL0[108] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5728 VSS WL0[108] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5729 VSS WL0[108] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5730 VSS WL0[108] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5731 VSS WL0[108] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5732 VSS WL0[108] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5733 VSS WL0[108] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5734 VSS WL0[108] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5735 VSS WL0[108] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5736 VSS WL0[108] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5737 VSS WL0[108] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5738 VSS WL0[108] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5739 VSS WL0[108] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5740 VSS WL0[108] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5741 VSS WL0[108] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5742 VSS WL0[108] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5743 VSS WL0[108] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5744 VSS WL0[108] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5745 VSS WL0[108] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5746 VSS WL0[108] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5747 VSS WL0[108] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5748 VSS WL0[108] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5749 VSS WL0[108] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5750 VSS WL0[108] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5751 VSS WL0[108] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5752 VSS WL0[108] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5753 VSS WL0[108] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5754 VSS WL0[108] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5755 VSS WL0[108] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5756 VSS WL0[108] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5757 VSS WL0[108] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5758 VSS WL0[108] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5759 VSS WL0[108] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5760 VSS WL0[108] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5761 VSS WL0[108] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5762 VSS WL0[108] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5763 VSS WL0[108] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5764 VSS WL0[108] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5765 VSS WL0[108] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5766 VSS WL0[108] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x6d0
XM5767 VSS WL0[109] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5768 VSS WL0[109] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5769 VSS WL0[109] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5770 VSS WL0[109] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5771 VSS WL0[109] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5772 VSS WL0[109] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5773 VSS WL0[109] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5774 VSS WL0[109] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5775 VSS WL0[109] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5776 VSS WL0[109] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5777 VSS WL0[109] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5778 VSS WL0[109] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5779 VSS WL0[109] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5780 VSS WL0[109] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5781 VSS WL0[109] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5782 VSS WL0[109] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5783 VSS WL0[109] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5784 VSS WL0[109] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5785 VSS WL0[109] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5786 VSS WL0[109] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5787 VSS WL0[109] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5788 VSS WL0[109] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5789 VSS WL0[109] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5790 VSS WL0[109] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5791 VSS WL0[109] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5792 VSS WL0[109] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5793 VSS WL0[109] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5794 VSS WL0[109] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5795 VSS WL0[109] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5796 VSS WL0[109] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5797 VSS WL0[109] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5798 VSS WL0[109] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5799 VSS WL0[109] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5800 VSS WL0[109] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5801 VSS WL0[109] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5802 VSS WL0[109] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5803 VSS WL0[109] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5804 VSS WL0[109] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5805 VSS WL0[109] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5806 VSS WL0[109] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5807 VSS WL0[109] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5808 VSS WL0[109] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5809 VSS WL0[109] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5810 VSS WL0[109] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5811 VSS WL0[109] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5812 VSS WL0[109] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5813 VSS WL0[109] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5814 VSS WL0[109] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5815 VSS WL0[109] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5816 VSS WL0[109] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5817 VSS WL0[109] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5818 VSS WL0[109] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5819 VSS WL0[109] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x6e0
XM5820 VSS WL0[110] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5821 VSS WL0[110] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5822 VSS WL0[110] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5823 VSS WL0[110] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5824 VSS WL0[110] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5825 VSS WL0[110] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5826 VSS WL0[110] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5827 VSS WL0[110] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5828 VSS WL0[110] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5829 VSS WL0[110] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5830 VSS WL0[110] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5831 VSS WL0[110] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5832 VSS WL0[110] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5833 VSS WL0[110] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5834 VSS WL0[110] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5835 VSS WL0[110] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5836 VSS WL0[110] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5837 VSS WL0[110] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5838 VSS WL0[110] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5839 VSS WL0[110] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5840 VSS WL0[110] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5841 VSS WL0[110] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5842 VSS WL0[110] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5843 VSS WL0[110] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5844 VSS WL0[110] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5845 VSS WL0[110] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5846 VSS WL0[110] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5847 VSS WL0[110] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5848 VSS WL0[110] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5849 VSS WL0[110] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5850 VSS WL0[110] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5851 VSS WL0[110] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5852 VSS WL0[110] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5853 VSS WL0[110] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5854 VSS WL0[110] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5855 VSS WL0[110] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5856 VSS WL0[110] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5857 VSS WL0[110] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5858 VSS WL0[110] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5859 VSS WL0[110] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5860 VSS WL0[110] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5861 VSS WL0[110] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5862 VSS WL0[110] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5863 VSS WL0[110] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5864 VSS WL0[110] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5865 VSS WL0[110] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5866 VSS WL0[110] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5867 VSS WL0[110] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5868 VSS WL0[110] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5869 VSS WL0[110] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5870 VSS WL0[110] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5871 VSS WL0[110] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5872 VSS WL0[110] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5873 VSS WL0[110] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x6f0
XM5874 VSS WL0[111] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5875 VSS WL0[111] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5876 VSS WL0[111] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5877 VSS WL0[111] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5878 VSS WL0[111] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5879 VSS WL0[111] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5880 VSS WL0[111] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5881 VSS WL0[111] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5882 VSS WL0[111] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5883 VSS WL0[111] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5884 VSS WL0[111] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5885 VSS WL0[111] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5886 VSS WL0[111] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5887 VSS WL0[111] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5888 VSS WL0[111] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5889 VSS WL0[111] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5890 VSS WL0[111] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5891 VSS WL0[111] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5892 VSS WL0[111] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5893 VSS WL0[111] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5894 VSS WL0[111] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5895 VSS WL0[111] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5896 VSS WL0[111] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5897 VSS WL0[111] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5898 VSS WL0[111] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5899 VSS WL0[111] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5900 VSS WL0[111] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5901 VSS WL0[111] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5902 VSS WL0[111] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5903 VSS WL0[111] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5904 VSS WL0[111] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5905 VSS WL0[111] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5906 VSS WL0[111] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5907 VSS WL0[111] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5908 VSS WL0[111] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5909 VSS WL0[111] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5910 VSS WL0[111] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5911 VSS WL0[111] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5912 VSS WL0[111] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5913 VSS WL0[111] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5914 VSS WL0[111] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5915 VSS WL0[111] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5916 VSS WL0[111] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5917 VSS WL0[111] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5918 VSS WL0[111] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5919 VSS WL0[111] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5920 VSS WL0[111] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5921 VSS WL0[111] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5922 VSS WL0[111] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x700
XM5923 VSS WL0[112] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5924 VSS WL0[112] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5925 VSS WL0[112] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5926 VSS WL0[112] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5927 VSS WL0[112] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5928 VSS WL0[112] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5929 VSS WL0[112] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5930 VSS WL0[112] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5931 VSS WL0[112] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5932 VSS WL0[112] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5933 VSS WL0[112] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5934 VSS WL0[112] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5935 VSS WL0[112] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5936 VSS WL0[112] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5937 VSS WL0[112] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5938 VSS WL0[112] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5939 VSS WL0[112] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5940 VSS WL0[112] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5941 VSS WL0[112] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5942 VSS WL0[112] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5943 VSS WL0[112] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5944 VSS WL0[112] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5945 VSS WL0[112] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5946 VSS WL0[112] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5947 VSS WL0[112] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5948 VSS WL0[112] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5949 VSS WL0[112] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5950 VSS WL0[112] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5951 VSS WL0[112] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5952 VSS WL0[112] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5953 VSS WL0[112] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5954 VSS WL0[112] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5955 VSS WL0[112] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5956 VSS WL0[112] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5957 VSS WL0[112] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5958 VSS WL0[112] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5959 VSS WL0[112] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5960 VSS WL0[112] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5961 VSS WL0[112] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5962 VSS WL0[112] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5963 VSS WL0[112] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5964 VSS WL0[112] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5965 VSS WL0[112] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x710
XM5966 VSS WL0[113] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5967 VSS WL0[113] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5968 VSS WL0[113] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5969 VSS WL0[113] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5970 VSS WL0[113] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5971 VSS WL0[113] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5972 VSS WL0[113] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5973 VSS WL0[113] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5974 VSS WL0[113] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5975 VSS WL0[113] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5976 VSS WL0[113] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5977 VSS WL0[113] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5978 VSS WL0[113] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5979 VSS WL0[113] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5980 VSS WL0[113] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5981 VSS WL0[113] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5982 VSS WL0[113] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5983 VSS WL0[113] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5984 VSS WL0[113] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5985 VSS WL0[113] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5986 VSS WL0[113] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5987 VSS WL0[113] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5988 VSS WL0[113] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5989 VSS WL0[113] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5990 VSS WL0[113] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5991 VSS WL0[113] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5992 VSS WL0[113] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5993 VSS WL0[113] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5994 VSS WL0[113] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5995 VSS WL0[113] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5996 VSS WL0[113] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5997 VSS WL0[113] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5998 VSS WL0[113] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM5999 VSS WL0[113] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6000 VSS WL0[113] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6001 VSS WL0[113] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6002 VSS WL0[113] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6003 VSS WL0[113] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6004 VSS WL0[113] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6005 VSS WL0[113] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6006 VSS WL0[113] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6007 VSS WL0[113] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6008 VSS WL0[113] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6009 VSS WL0[113] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6010 VSS WL0[113] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6011 VSS WL0[113] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6012 VSS WL0[113] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6013 VSS WL0[113] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6014 VSS WL0[113] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6015 VSS WL0[113] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6016 VSS WL0[113] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6017 VSS WL0[113] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6018 VSS WL0[113] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6019 VSS WL0[113] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6020 VSS WL0[113] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x720
XM6021 VSS WL0[114] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6022 VSS WL0[114] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6023 VSS WL0[114] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6024 VSS WL0[114] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6025 VSS WL0[114] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6026 VSS WL0[114] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6027 VSS WL0[114] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6028 VSS WL0[114] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6029 VSS WL0[114] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6030 VSS WL0[114] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6031 VSS WL0[114] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6032 VSS WL0[114] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6033 VSS WL0[114] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6034 VSS WL0[114] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6035 VSS WL0[114] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6036 VSS WL0[114] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6037 VSS WL0[114] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6038 VSS WL0[114] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6039 VSS WL0[114] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6040 VSS WL0[114] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6041 VSS WL0[114] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6042 VSS WL0[114] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6043 VSS WL0[114] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6044 VSS WL0[114] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6045 VSS WL0[114] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6046 VSS WL0[114] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6047 VSS WL0[114] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6048 VSS WL0[114] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6049 VSS WL0[114] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6050 VSS WL0[114] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6051 VSS WL0[114] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6052 VSS WL0[114] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6053 VSS WL0[114] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6054 VSS WL0[114] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6055 VSS WL0[114] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6056 VSS WL0[114] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6057 VSS WL0[114] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6058 VSS WL0[114] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6059 VSS WL0[114] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6060 VSS WL0[114] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6061 VSS WL0[114] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6062 VSS WL0[114] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6063 VSS WL0[114] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6064 VSS WL0[114] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6065 VSS WL0[114] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6066 VSS WL0[114] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6067 VSS WL0[114] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6068 VSS WL0[114] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x730
XM6069 VSS WL0[115] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6070 VSS WL0[115] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6071 VSS WL0[115] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6072 VSS WL0[115] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6073 VSS WL0[115] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6074 VSS WL0[115] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6075 VSS WL0[115] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6076 VSS WL0[115] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6077 VSS WL0[115] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6078 VSS WL0[115] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6079 VSS WL0[115] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6080 VSS WL0[115] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6081 VSS WL0[115] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6082 VSS WL0[115] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6083 VSS WL0[115] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6084 VSS WL0[115] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6085 VSS WL0[115] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6086 VSS WL0[115] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6087 VSS WL0[115] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6088 VSS WL0[115] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6089 VSS WL0[115] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6090 VSS WL0[115] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6091 VSS WL0[115] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6092 VSS WL0[115] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6093 VSS WL0[115] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6094 VSS WL0[115] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6095 VSS WL0[115] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6096 VSS WL0[115] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6097 VSS WL0[115] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6098 VSS WL0[115] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6099 VSS WL0[115] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6100 VSS WL0[115] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6101 VSS WL0[115] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6102 VSS WL0[115] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6103 VSS WL0[115] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6104 VSS WL0[115] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6105 VSS WL0[115] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6106 VSS WL0[115] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6107 VSS WL0[115] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6108 VSS WL0[115] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6109 VSS WL0[115] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6110 VSS WL0[115] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6111 VSS WL0[115] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6112 VSS WL0[115] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6113 VSS WL0[115] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6114 VSS WL0[115] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6115 VSS WL0[115] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6116 VSS WL0[115] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6117 VSS WL0[115] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6118 VSS WL0[115] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6119 VSS WL0[115] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6120 VSS WL0[115] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6121 VSS WL0[115] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6122 VSS WL0[115] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6123 VSS WL0[115] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6124 VSS WL0[115] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6125 VSS WL0[115] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6126 VSS WL0[115] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x740
XM6127 VSS WL0[116] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6128 VSS WL0[116] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6129 VSS WL0[116] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6130 VSS WL0[116] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6131 VSS WL0[116] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6132 VSS WL0[116] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6133 VSS WL0[116] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6134 VSS WL0[116] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6135 VSS WL0[116] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6136 VSS WL0[116] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6137 VSS WL0[116] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6138 VSS WL0[116] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6139 VSS WL0[116] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6140 VSS WL0[116] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6141 VSS WL0[116] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6142 VSS WL0[116] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6143 VSS WL0[116] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6144 VSS WL0[116] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6145 VSS WL0[116] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6146 VSS WL0[116] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6147 VSS WL0[116] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6148 VSS WL0[116] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6149 VSS WL0[116] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6150 VSS WL0[116] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6151 VSS WL0[116] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6152 VSS WL0[116] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6153 VSS WL0[116] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6154 VSS WL0[116] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6155 VSS WL0[116] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6156 VSS WL0[116] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6157 VSS WL0[116] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6158 VSS WL0[116] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6159 VSS WL0[116] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6160 VSS WL0[116] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6161 VSS WL0[116] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6162 VSS WL0[116] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6163 VSS WL0[116] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6164 VSS WL0[116] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6165 VSS WL0[116] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6166 VSS WL0[116] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6167 VSS WL0[116] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6168 VSS WL0[116] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6169 VSS WL0[116] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6170 VSS WL0[116] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6171 VSS WL0[116] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6172 VSS WL0[116] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6173 VSS WL0[116] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6174 VSS WL0[116] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6175 VSS WL0[116] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6176 VSS WL0[116] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6177 VSS WL0[116] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6178 VSS WL0[116] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6179 VSS WL0[116] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6180 VSS WL0[116] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6181 VSS WL0[116] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6182 VSS WL0[116] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6183 VSS WL0[116] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x750
XM6184 VSS WL0[117] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6185 VSS WL0[117] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6186 VSS WL0[117] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6187 VSS WL0[117] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6188 VSS WL0[117] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6189 VSS WL0[117] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6190 VSS WL0[117] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6191 VSS WL0[117] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6192 VSS WL0[117] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6193 VSS WL0[117] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6194 VSS WL0[117] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6195 VSS WL0[117] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6196 VSS WL0[117] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6197 VSS WL0[117] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6198 VSS WL0[117] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6199 VSS WL0[117] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6200 VSS WL0[117] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6201 VSS WL0[117] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6202 VSS WL0[117] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6203 VSS WL0[117] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6204 VSS WL0[117] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6205 VSS WL0[117] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6206 VSS WL0[117] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6207 VSS WL0[117] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6208 VSS WL0[117] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6209 VSS WL0[117] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6210 VSS WL0[117] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6211 VSS WL0[117] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6212 VSS WL0[117] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6213 VSS WL0[117] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6214 VSS WL0[117] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6215 VSS WL0[117] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6216 VSS WL0[117] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6217 VSS WL0[117] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6218 VSS WL0[117] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6219 VSS WL0[117] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6220 VSS WL0[117] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6221 VSS WL0[117] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6222 VSS WL0[117] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6223 VSS WL0[117] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6224 VSS WL0[117] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6225 VSS WL0[117] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6226 VSS WL0[117] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6227 VSS WL0[117] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6228 VSS WL0[117] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6229 VSS WL0[117] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6230 VSS WL0[117] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6231 VSS WL0[117] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6232 VSS WL0[117] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6233 VSS WL0[117] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6234 VSS WL0[117] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6235 VSS WL0[117] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6236 VSS WL0[117] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6237 VSS WL0[117] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6238 VSS WL0[117] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6239 VSS WL0[117] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6240 VSS WL0[117] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6241 VSS WL0[117] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6242 VSS WL0[117] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6243 VSS WL0[117] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6244 VSS WL0[117] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6245 VSS WL0[117] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x760
XM6246 VSS WL0[118] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6247 VSS WL0[118] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6248 VSS WL0[118] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6249 VSS WL0[118] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6250 VSS WL0[118] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6251 VSS WL0[118] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6252 VSS WL0[118] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6253 VSS WL0[118] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6254 VSS WL0[118] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6255 VSS WL0[118] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6256 VSS WL0[118] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6257 VSS WL0[118] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6258 VSS WL0[118] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6259 VSS WL0[118] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6260 VSS WL0[118] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6261 VSS WL0[118] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6262 VSS WL0[118] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6263 VSS WL0[118] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6264 VSS WL0[118] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6265 VSS WL0[118] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6266 VSS WL0[118] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6267 VSS WL0[118] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6268 VSS WL0[118] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6269 VSS WL0[118] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6270 VSS WL0[118] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6271 VSS WL0[118] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6272 VSS WL0[118] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6273 VSS WL0[118] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6274 VSS WL0[118] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6275 VSS WL0[118] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6276 VSS WL0[118] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6277 VSS WL0[118] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6278 VSS WL0[118] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6279 VSS WL0[118] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6280 VSS WL0[118] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6281 VSS WL0[118] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6282 VSS WL0[118] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6283 VSS WL0[118] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6284 VSS WL0[118] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6285 VSS WL0[118] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6286 VSS WL0[118] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6287 VSS WL0[118] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6288 VSS WL0[118] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6289 VSS WL0[118] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6290 VSS WL0[118] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6291 VSS WL0[118] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6292 VSS WL0[118] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6293 VSS WL0[118] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6294 VSS WL0[118] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6295 VSS WL0[118] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6296 VSS WL0[118] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6297 VSS WL0[118] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6298 VSS WL0[118] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6299 VSS WL0[118] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6300 VSS WL0[118] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x770
XM6301 VSS WL0[119] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6302 VSS WL0[119] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6303 VSS WL0[119] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6304 VSS WL0[119] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6305 VSS WL0[119] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6306 VSS WL0[119] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6307 VSS WL0[119] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6308 VSS WL0[119] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6309 VSS WL0[119] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6310 VSS WL0[119] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6311 VSS WL0[119] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6312 VSS WL0[119] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6313 VSS WL0[119] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6314 VSS WL0[119] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6315 VSS WL0[119] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6316 VSS WL0[119] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6317 VSS WL0[119] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6318 VSS WL0[119] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6319 VSS WL0[119] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6320 VSS WL0[119] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6321 VSS WL0[119] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6322 VSS WL0[119] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6323 VSS WL0[119] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6324 VSS WL0[119] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6325 VSS WL0[119] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6326 VSS WL0[119] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6327 VSS WL0[119] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6328 VSS WL0[119] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6329 VSS WL0[119] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6330 VSS WL0[119] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6331 VSS WL0[119] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6332 VSS WL0[119] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6333 VSS WL0[119] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6334 VSS WL0[119] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6335 VSS WL0[119] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6336 VSS WL0[119] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6337 VSS WL0[119] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6338 VSS WL0[119] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6339 VSS WL0[119] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6340 VSS WL0[119] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6341 VSS WL0[119] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6342 VSS WL0[119] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6343 VSS WL0[119] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6344 VSS WL0[119] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6345 VSS WL0[119] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6346 VSS WL0[119] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6347 VSS WL0[119] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6348 VSS WL0[119] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6349 VSS WL0[119] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6350 VSS WL0[119] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6351 VSS WL0[119] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6352 VSS WL0[119] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6353 VSS WL0[119] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6354 VSS WL0[119] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x780
XM6355 VSS WL0[120] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6356 VSS WL0[120] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6357 VSS WL0[120] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6358 VSS WL0[120] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6359 VSS WL0[120] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6360 VSS WL0[120] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6361 VSS WL0[120] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6362 VSS WL0[120] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6363 VSS WL0[120] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6364 VSS WL0[120] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6365 VSS WL0[120] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6366 VSS WL0[120] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6367 VSS WL0[120] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6368 VSS WL0[120] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6369 VSS WL0[120] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6370 VSS WL0[120] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6371 VSS WL0[120] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6372 VSS WL0[120] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6373 VSS WL0[120] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6374 VSS WL0[120] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6375 VSS WL0[120] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6376 VSS WL0[120] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6377 VSS WL0[120] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6378 VSS WL0[120] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6379 VSS WL0[120] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6380 VSS WL0[120] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6381 VSS WL0[120] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6382 VSS WL0[120] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6383 VSS WL0[120] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6384 VSS WL0[120] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6385 VSS WL0[120] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6386 VSS WL0[120] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6387 VSS WL0[120] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6388 VSS WL0[120] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6389 VSS WL0[120] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6390 VSS WL0[120] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6391 VSS WL0[120] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6392 VSS WL0[120] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6393 VSS WL0[120] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6394 VSS WL0[120] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6395 VSS WL0[120] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6396 VSS WL0[120] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6397 VSS WL0[120] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6398 VSS WL0[120] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6399 VSS WL0[120] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6400 VSS WL0[120] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6401 VSS WL0[120] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6402 VSS WL0[120] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6403 VSS WL0[120] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6404 VSS WL0[120] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6405 VSS WL0[120] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6406 VSS WL0[120] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6407 VSS WL0[120] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6408 VSS WL0[120] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6409 VSS WL0[120] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6410 VSS WL0[120] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6411 VSS WL0[120] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6412 VSS WL0[120] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6413 VSS WL0[120] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6414 VSS WL0[120] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6415 VSS WL0[120] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x790
XM6416 VSS WL0[121] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6417 VSS WL0[121] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6418 VSS WL0[121] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6419 VSS WL0[121] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6420 VSS WL0[121] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6421 VSS WL0[121] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6422 VSS WL0[121] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6423 VSS WL0[121] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6424 VSS WL0[121] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6425 VSS WL0[121] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6426 VSS WL0[121] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6427 VSS WL0[121] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6428 VSS WL0[121] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6429 VSS WL0[121] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6430 VSS WL0[121] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6431 VSS WL0[121] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6432 VSS WL0[121] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6433 VSS WL0[121] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6434 VSS WL0[121] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6435 VSS WL0[121] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6436 VSS WL0[121] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6437 VSS WL0[121] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6438 VSS WL0[121] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6439 VSS WL0[121] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6440 VSS WL0[121] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6441 VSS WL0[121] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6442 VSS WL0[121] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6443 VSS WL0[121] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6444 VSS WL0[121] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6445 VSS WL0[121] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6446 VSS WL0[121] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6447 VSS WL0[121] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6448 VSS WL0[121] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6449 VSS WL0[121] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6450 VSS WL0[121] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6451 VSS WL0[121] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6452 VSS WL0[121] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6453 VSS WL0[121] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6454 VSS WL0[121] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6455 VSS WL0[121] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6456 VSS WL0[121] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6457 VSS WL0[121] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6458 VSS WL0[121] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6459 VSS WL0[121] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6460 VSS WL0[121] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6461 VSS WL0[121] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6462 VSS WL0[121] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6463 VSS WL0[121] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6464 VSS WL0[121] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6465 VSS WL0[121] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6466 VSS WL0[121] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6467 VSS WL0[121] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6468 VSS WL0[121] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6469 VSS WL0[121] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6470 VSS WL0[121] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6471 VSS WL0[121] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6472 VSS WL0[121] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6473 VSS WL0[121] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6474 VSS WL0[121] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6475 VSS WL0[121] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6476 VSS WL0[121] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x7a0
XM6477 VSS WL0[122] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6478 VSS WL0[122] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6479 VSS WL0[122] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6480 VSS WL0[122] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6481 VSS WL0[122] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6482 VSS WL0[122] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6483 VSS WL0[122] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6484 VSS WL0[122] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6485 VSS WL0[122] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6486 VSS WL0[122] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6487 VSS WL0[122] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6488 VSS WL0[122] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6489 VSS WL0[122] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6490 VSS WL0[122] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6491 VSS WL0[122] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6492 VSS WL0[122] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6493 VSS WL0[122] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6494 VSS WL0[122] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6495 VSS WL0[122] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6496 VSS WL0[122] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6497 VSS WL0[122] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6498 VSS WL0[122] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6499 VSS WL0[122] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6500 VSS WL0[122] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6501 VSS WL0[122] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6502 VSS WL0[122] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6503 VSS WL0[122] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6504 VSS WL0[122] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6505 VSS WL0[122] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6506 VSS WL0[122] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6507 VSS WL0[122] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6508 VSS WL0[122] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6509 VSS WL0[122] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6510 VSS WL0[122] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6511 VSS WL0[122] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6512 VSS WL0[122] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6513 VSS WL0[122] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6514 VSS WL0[122] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6515 VSS WL0[122] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6516 VSS WL0[122] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6517 VSS WL0[122] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6518 VSS WL0[122] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6519 VSS WL0[122] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6520 VSS WL0[122] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6521 VSS WL0[122] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6522 VSS WL0[122] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6523 VSS WL0[122] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6524 VSS WL0[122] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6525 VSS WL0[122] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6526 VSS WL0[122] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6527 VSS WL0[122] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6528 VSS WL0[122] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6529 VSS WL0[122] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6530 VSS WL0[122] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6531 VSS WL0[122] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6532 VSS WL0[122] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6533 VSS WL0[122] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6534 VSS WL0[122] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6535 VSS WL0[122] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6536 VSS WL0[122] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x7b0
XM6537 VSS WL0[123] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6538 VSS WL0[123] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6539 VSS WL0[123] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6540 VSS WL0[123] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6541 VSS WL0[123] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6542 VSS WL0[123] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6543 VSS WL0[123] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6544 VSS WL0[123] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6545 VSS WL0[123] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6546 VSS WL0[123] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6547 VSS WL0[123] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6548 VSS WL0[123] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6549 VSS WL0[123] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6550 VSS WL0[123] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6551 VSS WL0[123] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6552 VSS WL0[123] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6553 VSS WL0[123] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6554 VSS WL0[123] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6555 VSS WL0[123] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6556 VSS WL0[123] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6557 VSS WL0[123] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6558 VSS WL0[123] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6559 VSS WL0[123] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6560 VSS WL0[123] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6561 VSS WL0[123] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6562 VSS WL0[123] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6563 VSS WL0[123] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6564 VSS WL0[123] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6565 VSS WL0[123] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6566 VSS WL0[123] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6567 VSS WL0[123] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6568 VSS WL0[123] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6569 VSS WL0[123] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6570 VSS WL0[123] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6571 VSS WL0[123] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6572 VSS WL0[123] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6573 VSS WL0[123] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6574 VSS WL0[123] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6575 VSS WL0[123] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6576 VSS WL0[123] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6577 VSS WL0[123] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6578 VSS WL0[123] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6579 VSS WL0[123] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6580 VSS WL0[123] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6581 VSS WL0[123] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6582 VSS WL0[123] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6583 VSS WL0[123] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6584 VSS WL0[123] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6585 VSS WL0[123] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6586 VSS WL0[123] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6587 VSS WL0[123] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6588 VSS WL0[123] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6589 VSS WL0[123] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6590 VSS WL0[123] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6591 VSS WL0[123] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6592 VSS WL0[123] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6593 VSS WL0[123] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6594 VSS WL0[123] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6595 VSS WL0[123] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6596 VSS WL0[123] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6597 VSS WL0[123] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6598 VSS WL0[123] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6599 VSS WL0[123] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x7c0
XM6600 VSS WL0[124] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6601 VSS WL0[124] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6602 VSS WL0[124] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6603 VSS WL0[124] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6604 VSS WL0[124] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6605 VSS WL0[124] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6606 VSS WL0[124] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6607 VSS WL0[124] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6608 VSS WL0[124] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6609 VSS WL0[124] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6610 VSS WL0[124] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6611 VSS WL0[124] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6612 VSS WL0[124] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6613 VSS WL0[124] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6614 VSS WL0[124] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6615 VSS WL0[124] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6616 VSS WL0[124] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6617 VSS WL0[124] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6618 VSS WL0[124] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6619 VSS WL0[124] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6620 VSS WL0[124] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6621 VSS WL0[124] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6622 VSS WL0[124] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6623 VSS WL0[124] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6624 VSS WL0[124] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6625 VSS WL0[124] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6626 VSS WL0[124] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6627 VSS WL0[124] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6628 VSS WL0[124] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6629 VSS WL0[124] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6630 VSS WL0[124] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6631 VSS WL0[124] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6632 VSS WL0[124] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6633 VSS WL0[124] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6634 VSS WL0[124] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6635 VSS WL0[124] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6636 VSS WL0[124] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6637 VSS WL0[124] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6638 VSS WL0[124] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6639 VSS WL0[124] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6640 VSS WL0[124] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6641 VSS WL0[124] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6642 VSS WL0[124] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6643 VSS WL0[124] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6644 VSS WL0[124] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6645 VSS WL0[124] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6646 VSS WL0[124] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6647 VSS WL0[124] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6648 VSS WL0[124] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6649 VSS WL0[124] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6650 VSS WL0[124] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6651 VSS WL0[124] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6652 VSS WL0[124] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6653 VSS WL0[124] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6654 VSS WL0[124] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6655 VSS WL0[124] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6656 VSS WL0[124] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6657 VSS WL0[124] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6658 VSS WL0[124] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6659 VSS WL0[124] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6660 VSS WL0[124] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6661 VSS WL0[124] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x7d0
XM6662 VSS WL0[125] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6663 VSS WL0[125] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6664 VSS WL0[125] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6665 VSS WL0[125] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6666 VSS WL0[125] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6667 VSS WL0[125] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6668 VSS WL0[125] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6669 VSS WL0[125] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6670 VSS WL0[125] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6671 VSS WL0[125] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6672 VSS WL0[125] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6673 VSS WL0[125] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6674 VSS WL0[125] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6675 VSS WL0[125] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6676 VSS WL0[125] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6677 VSS WL0[125] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6678 VSS WL0[125] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6679 VSS WL0[125] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6680 VSS WL0[125] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6681 VSS WL0[125] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6682 VSS WL0[125] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6683 VSS WL0[125] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6684 VSS WL0[125] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6685 VSS WL0[125] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6686 VSS WL0[125] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6687 VSS WL0[125] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6688 VSS WL0[125] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6689 VSS WL0[125] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6690 VSS WL0[125] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6691 VSS WL0[125] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6692 VSS WL0[125] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6693 VSS WL0[125] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6694 VSS WL0[125] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6695 VSS WL0[125] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6696 VSS WL0[125] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6697 VSS WL0[125] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6698 VSS WL0[125] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6699 VSS WL0[125] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6700 VSS WL0[125] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6701 VSS WL0[125] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6702 VSS WL0[125] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6703 VSS WL0[125] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6704 VSS WL0[125] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6705 VSS WL0[125] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6706 VSS WL0[125] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6707 VSS WL0[125] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6708 VSS WL0[125] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6709 VSS WL0[125] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6710 VSS WL0[125] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6711 VSS WL0[125] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6712 VSS WL0[125] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6713 VSS WL0[125] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6714 VSS WL0[125] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6715 VSS WL0[125] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6716 VSS WL0[125] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6717 VSS WL0[125] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6718 VSS WL0[125] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6719 VSS WL0[125] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6720 VSS WL0[125] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x7e0
XM6721 VSS WL0[126] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6722 VSS WL0[126] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6723 VSS WL0[126] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6724 VSS WL0[126] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6725 VSS WL0[126] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6726 VSS WL0[126] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6727 VSS WL0[126] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6728 VSS WL0[126] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6729 VSS WL0[126] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6730 VSS WL0[126] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6731 VSS WL0[126] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6732 VSS WL0[126] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6733 VSS WL0[126] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6734 VSS WL0[126] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6735 VSS WL0[126] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6736 VSS WL0[126] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6737 VSS WL0[126] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6738 VSS WL0[126] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6739 VSS WL0[126] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6740 VSS WL0[126] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6741 VSS WL0[126] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6742 VSS WL0[126] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6743 VSS WL0[126] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6744 VSS WL0[126] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6745 VSS WL0[126] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6746 VSS WL0[126] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6747 VSS WL0[126] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6748 VSS WL0[126] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6749 VSS WL0[126] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6750 VSS WL0[126] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6751 VSS WL0[126] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6752 VSS WL0[126] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6753 VSS WL0[126] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6754 VSS WL0[126] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6755 VSS WL0[126] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6756 VSS WL0[126] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6757 VSS WL0[126] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6758 VSS WL0[126] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6759 VSS WL0[126] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6760 VSS WL0[126] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6761 VSS WL0[126] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6762 VSS WL0[126] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6763 VSS WL0[126] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6764 VSS WL0[126] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6765 VSS WL0[126] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6766 VSS WL0[126] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6767 VSS WL0[126] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6768 VSS WL0[126] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6769 VSS WL0[126] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6770 VSS WL0[126] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6771 VSS WL0[126] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6772 VSS WL0[126] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6773 VSS WL0[126] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6774 VSS WL0[126] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x7f0
XM6775 VSS WL0[127] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6776 VSS WL0[127] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6777 VSS WL0[127] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6778 VSS WL0[127] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6779 VSS WL0[127] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6780 VSS WL0[127] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6781 VSS WL0[127] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6782 VSS WL0[127] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6783 VSS WL0[127] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6784 VSS WL0[127] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6785 VSS WL0[127] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6786 VSS WL0[127] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6787 VSS WL0[127] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6788 VSS WL0[127] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6789 VSS WL0[127] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6790 VSS WL0[127] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6791 VSS WL0[127] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6792 VSS WL0[127] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6793 VSS WL0[127] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6794 VSS WL0[127] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6795 VSS WL0[127] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6796 VSS WL0[127] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6797 VSS WL0[127] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6798 VSS WL0[127] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6799 VSS WL0[127] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6800 VSS WL0[127] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6801 VSS WL0[127] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6802 VSS WL0[127] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6803 VSS WL0[127] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6804 VSS WL0[127] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6805 VSS WL0[127] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6806 VSS WL0[127] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6807 VSS WL0[127] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6808 VSS WL0[127] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6809 VSS WL0[127] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6810 VSS WL0[127] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6811 VSS WL0[127] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6812 VSS WL0[127] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6813 VSS WL0[127] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6814 VSS WL0[127] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6815 VSS WL0[127] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6816 VSS WL0[127] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6817 VSS WL0[127] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6818 VSS WL0[127] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6819 VSS WL0[127] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6820 VSS WL0[127] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6821 VSS WL0[127] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6822 VSS WL0[127] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6823 VSS WL0[127] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6824 VSS WL0[127] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6825 VSS WL0[127] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6826 VSS WL0[127] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6827 VSS WL0[127] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6828 VSS WL0[127] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6829 VSS WL0[127] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6830 VSS WL0[127] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6831 VSS WL0[127] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6832 VSS WL0[127] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6833 VSS WL0[127] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x800
XM6834 VSS WL0[128] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6835 VSS WL0[128] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6836 VSS WL0[128] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6837 VSS WL0[128] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6838 VSS WL0[128] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6839 VSS WL0[128] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6840 VSS WL0[128] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6841 VSS WL0[128] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6842 VSS WL0[128] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6843 VSS WL0[128] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6844 VSS WL0[128] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6845 VSS WL0[128] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6846 VSS WL0[128] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6847 VSS WL0[128] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6848 VSS WL0[128] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6849 VSS WL0[128] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6850 VSS WL0[128] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6851 VSS WL0[128] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6852 VSS WL0[128] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6853 VSS WL0[128] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6854 VSS WL0[128] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6855 VSS WL0[128] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6856 VSS WL0[128] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6857 VSS WL0[128] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6858 VSS WL0[128] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6859 VSS WL0[128] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6860 VSS WL0[128] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6861 VSS WL0[128] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6862 VSS WL0[128] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6863 VSS WL0[128] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6864 VSS WL0[128] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6865 VSS WL0[128] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6866 VSS WL0[128] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6867 VSS WL0[128] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6868 VSS WL0[128] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6869 VSS WL0[128] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6870 VSS WL0[128] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6871 VSS WL0[128] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6872 VSS WL0[128] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6873 VSS WL0[128] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6874 VSS WL0[128] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6875 VSS WL0[128] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6876 VSS WL0[128] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6877 VSS WL0[128] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6878 VSS WL0[128] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6879 VSS WL0[128] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6880 VSS WL0[128] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6881 VSS WL0[128] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6882 VSS WL0[128] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6883 VSS WL0[128] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6884 VSS WL0[128] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6885 VSS WL0[128] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6886 VSS WL0[128] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6887 VSS WL0[128] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6888 VSS WL0[128] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x810
XM6889 VSS WL0[129] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6890 VSS WL0[129] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6891 VSS WL0[129] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6892 VSS WL0[129] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6893 VSS WL0[129] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6894 VSS WL0[129] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6895 VSS WL0[129] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6896 VSS WL0[129] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6897 VSS WL0[129] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6898 VSS WL0[129] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6899 VSS WL0[129] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6900 VSS WL0[129] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6901 VSS WL0[129] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6902 VSS WL0[129] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6903 VSS WL0[129] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6904 VSS WL0[129] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6905 VSS WL0[129] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6906 VSS WL0[129] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6907 VSS WL0[129] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6908 VSS WL0[129] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6909 VSS WL0[129] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6910 VSS WL0[129] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6911 VSS WL0[129] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6912 VSS WL0[129] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6913 VSS WL0[129] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6914 VSS WL0[129] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6915 VSS WL0[129] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6916 VSS WL0[129] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6917 VSS WL0[129] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6918 VSS WL0[129] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6919 VSS WL0[129] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6920 VSS WL0[129] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6921 VSS WL0[129] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6922 VSS WL0[129] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6923 VSS WL0[129] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6924 VSS WL0[129] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6925 VSS WL0[129] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6926 VSS WL0[129] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6927 VSS WL0[129] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6928 VSS WL0[129] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6929 VSS WL0[129] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6930 VSS WL0[129] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6931 VSS WL0[129] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6932 VSS WL0[129] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6933 VSS WL0[129] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6934 VSS WL0[129] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6935 VSS WL0[129] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6936 VSS WL0[129] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6937 VSS WL0[129] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6938 VSS WL0[129] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6939 VSS WL0[129] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6940 VSS WL0[129] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6941 VSS WL0[129] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6942 VSS WL0[129] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6943 VSS WL0[129] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6944 VSS WL0[129] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6945 VSS WL0[129] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6946 VSS WL0[129] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6947 VSS WL0[129] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6948 VSS WL0[129] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6949 VSS WL0[129] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6950 VSS WL0[129] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6951 VSS WL0[129] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x820
XM6952 VSS WL0[130] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6953 VSS WL0[130] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6954 VSS WL0[130] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6955 VSS WL0[130] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6956 VSS WL0[130] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6957 VSS WL0[130] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6958 VSS WL0[130] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6959 VSS WL0[130] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6960 VSS WL0[130] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6961 VSS WL0[130] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6962 VSS WL0[130] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6963 VSS WL0[130] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6964 VSS WL0[130] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6965 VSS WL0[130] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6966 VSS WL0[130] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6967 VSS WL0[130] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6968 VSS WL0[130] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6969 VSS WL0[130] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6970 VSS WL0[130] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6971 VSS WL0[130] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6972 VSS WL0[130] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6973 VSS WL0[130] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6974 VSS WL0[130] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6975 VSS WL0[130] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6976 VSS WL0[130] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6977 VSS WL0[130] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6978 VSS WL0[130] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6979 VSS WL0[130] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6980 VSS WL0[130] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6981 VSS WL0[130] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6982 VSS WL0[130] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6983 VSS WL0[130] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6984 VSS WL0[130] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6985 VSS WL0[130] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6986 VSS WL0[130] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6987 VSS WL0[130] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6988 VSS WL0[130] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6989 VSS WL0[130] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6990 VSS WL0[130] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6991 VSS WL0[130] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6992 VSS WL0[130] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6993 VSS WL0[130] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6994 VSS WL0[130] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6995 VSS WL0[130] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6996 VSS WL0[130] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6997 VSS WL0[130] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6998 VSS WL0[130] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM6999 VSS WL0[130] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7000 VSS WL0[130] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7001 VSS WL0[130] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7002 VSS WL0[130] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7003 VSS WL0[130] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7004 VSS WL0[130] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x830
XM7005 VSS WL0[131] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7006 VSS WL0[131] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7007 VSS WL0[131] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7008 VSS WL0[131] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7009 VSS WL0[131] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7010 VSS WL0[131] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7011 VSS WL0[131] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7012 VSS WL0[131] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7013 VSS WL0[131] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7014 VSS WL0[131] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7015 VSS WL0[131] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7016 VSS WL0[131] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7017 VSS WL0[131] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7018 VSS WL0[131] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7019 VSS WL0[131] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7020 VSS WL0[131] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7021 VSS WL0[131] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7022 VSS WL0[131] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7023 VSS WL0[131] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7024 VSS WL0[131] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7025 VSS WL0[131] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7026 VSS WL0[131] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7027 VSS WL0[131] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7028 VSS WL0[131] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7029 VSS WL0[131] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7030 VSS WL0[131] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7031 VSS WL0[131] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7032 VSS WL0[131] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7033 VSS WL0[131] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7034 VSS WL0[131] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7035 VSS WL0[131] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7036 VSS WL0[131] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7037 VSS WL0[131] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7038 VSS WL0[131] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7039 VSS WL0[131] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7040 VSS WL0[131] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7041 VSS WL0[131] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7042 VSS WL0[131] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7043 VSS WL0[131] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7044 VSS WL0[131] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7045 VSS WL0[131] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7046 VSS WL0[131] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7047 VSS WL0[131] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7048 VSS WL0[131] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7049 VSS WL0[131] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7050 VSS WL0[131] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7051 VSS WL0[131] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7052 VSS WL0[131] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7053 VSS WL0[131] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x840
XM7054 VSS WL0[132] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7055 VSS WL0[132] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7056 VSS WL0[132] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7057 VSS WL0[132] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7058 VSS WL0[132] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7059 VSS WL0[132] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7060 VSS WL0[132] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7061 VSS WL0[132] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7062 VSS WL0[132] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7063 VSS WL0[132] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7064 VSS WL0[132] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7065 VSS WL0[132] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7066 VSS WL0[132] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7067 VSS WL0[132] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7068 VSS WL0[132] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7069 VSS WL0[132] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7070 VSS WL0[132] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7071 VSS WL0[132] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7072 VSS WL0[132] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7073 VSS WL0[132] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7074 VSS WL0[132] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7075 VSS WL0[132] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7076 VSS WL0[132] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7077 VSS WL0[132] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7078 VSS WL0[132] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7079 VSS WL0[132] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7080 VSS WL0[132] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7081 VSS WL0[132] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7082 VSS WL0[132] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7083 VSS WL0[132] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7084 VSS WL0[132] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7085 VSS WL0[132] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7086 VSS WL0[132] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7087 VSS WL0[132] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7088 VSS WL0[132] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7089 VSS WL0[132] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7090 VSS WL0[132] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7091 VSS WL0[132] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7092 VSS WL0[132] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7093 VSS WL0[132] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7094 VSS WL0[132] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7095 VSS WL0[132] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7096 VSS WL0[132] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7097 VSS WL0[132] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7098 VSS WL0[132] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7099 VSS WL0[132] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7100 VSS WL0[132] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7101 VSS WL0[132] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7102 VSS WL0[132] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7103 VSS WL0[132] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7104 VSS WL0[132] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7105 VSS WL0[132] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7106 VSS WL0[132] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7107 VSS WL0[132] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7108 VSS WL0[132] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7109 VSS WL0[132] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x850
XM7110 VSS WL0[133] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7111 VSS WL0[133] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7112 VSS WL0[133] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7113 VSS WL0[133] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7114 VSS WL0[133] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7115 VSS WL0[133] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7116 VSS WL0[133] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7117 VSS WL0[133] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7118 VSS WL0[133] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7119 VSS WL0[133] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7120 VSS WL0[133] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7121 VSS WL0[133] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7122 VSS WL0[133] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7123 VSS WL0[133] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7124 VSS WL0[133] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7125 VSS WL0[133] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7126 VSS WL0[133] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7127 VSS WL0[133] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7128 VSS WL0[133] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7129 VSS WL0[133] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7130 VSS WL0[133] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7131 VSS WL0[133] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7132 VSS WL0[133] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7133 VSS WL0[133] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7134 VSS WL0[133] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7135 VSS WL0[133] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7136 VSS WL0[133] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7137 VSS WL0[133] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7138 VSS WL0[133] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7139 VSS WL0[133] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7140 VSS WL0[133] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7141 VSS WL0[133] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7142 VSS WL0[133] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7143 VSS WL0[133] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7144 VSS WL0[133] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7145 VSS WL0[133] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7146 VSS WL0[133] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7147 VSS WL0[133] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7148 VSS WL0[133] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7149 VSS WL0[133] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7150 VSS WL0[133] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7151 VSS WL0[133] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7152 VSS WL0[133] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7153 VSS WL0[133] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7154 VSS WL0[133] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7155 VSS WL0[133] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7156 VSS WL0[133] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x860
XM7157 VSS WL0[134] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7158 VSS WL0[134] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7159 VSS WL0[134] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7160 VSS WL0[134] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7161 VSS WL0[134] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7162 VSS WL0[134] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7163 VSS WL0[134] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7164 VSS WL0[134] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7165 VSS WL0[134] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7166 VSS WL0[134] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7167 VSS WL0[134] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7168 VSS WL0[134] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7169 VSS WL0[134] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7170 VSS WL0[134] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7171 VSS WL0[134] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7172 VSS WL0[134] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7173 VSS WL0[134] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7174 VSS WL0[134] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7175 VSS WL0[134] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7176 VSS WL0[134] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7177 VSS WL0[134] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7178 VSS WL0[134] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7179 VSS WL0[134] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7180 VSS WL0[134] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7181 VSS WL0[134] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7182 VSS WL0[134] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7183 VSS WL0[134] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7184 VSS WL0[134] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7185 VSS WL0[134] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7186 VSS WL0[134] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7187 VSS WL0[134] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7188 VSS WL0[134] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7189 VSS WL0[134] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7190 VSS WL0[134] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7191 VSS WL0[134] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7192 VSS WL0[134] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7193 VSS WL0[134] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7194 VSS WL0[134] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7195 VSS WL0[134] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7196 VSS WL0[134] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7197 VSS WL0[134] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7198 VSS WL0[134] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7199 VSS WL0[134] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7200 VSS WL0[134] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7201 VSS WL0[134] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x870
XM7202 VSS WL0[135] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7203 VSS WL0[135] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7204 VSS WL0[135] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7205 VSS WL0[135] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7206 VSS WL0[135] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7207 VSS WL0[135] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7208 VSS WL0[135] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7209 VSS WL0[135] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7210 VSS WL0[135] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7211 VSS WL0[135] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7212 VSS WL0[135] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7213 VSS WL0[135] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7214 VSS WL0[135] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7215 VSS WL0[135] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7216 VSS WL0[135] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7217 VSS WL0[135] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7218 VSS WL0[135] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7219 VSS WL0[135] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7220 VSS WL0[135] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7221 VSS WL0[135] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7222 VSS WL0[135] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7223 VSS WL0[135] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7224 VSS WL0[135] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7225 VSS WL0[135] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7226 VSS WL0[135] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7227 VSS WL0[135] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7228 VSS WL0[135] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7229 VSS WL0[135] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7230 VSS WL0[135] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7231 VSS WL0[135] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7232 VSS WL0[135] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7233 VSS WL0[135] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7234 VSS WL0[135] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7235 VSS WL0[135] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7236 VSS WL0[135] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7237 VSS WL0[135] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7238 VSS WL0[135] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7239 VSS WL0[135] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7240 VSS WL0[135] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7241 VSS WL0[135] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7242 VSS WL0[135] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7243 VSS WL0[135] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7244 VSS WL0[135] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7245 VSS WL0[135] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7246 VSS WL0[135] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7247 VSS WL0[135] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7248 VSS WL0[135] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7249 VSS WL0[135] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7250 VSS WL0[135] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7251 VSS WL0[135] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7252 VSS WL0[135] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7253 VSS WL0[135] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7254 VSS WL0[135] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7255 VSS WL0[135] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7256 VSS WL0[135] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7257 VSS WL0[135] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7258 VSS WL0[135] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7259 VSS WL0[135] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x880
XM7260 VSS WL0[136] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7261 VSS WL0[136] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7262 VSS WL0[136] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7263 VSS WL0[136] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7264 VSS WL0[136] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7265 VSS WL0[136] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7266 VSS WL0[136] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7267 VSS WL0[136] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7268 VSS WL0[136] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7269 VSS WL0[136] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7270 VSS WL0[136] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7271 VSS WL0[136] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7272 VSS WL0[136] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7273 VSS WL0[136] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7274 VSS WL0[136] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7275 VSS WL0[136] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7276 VSS WL0[136] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7277 VSS WL0[136] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7278 VSS WL0[136] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7279 VSS WL0[136] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7280 VSS WL0[136] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7281 VSS WL0[136] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7282 VSS WL0[136] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7283 VSS WL0[136] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7284 VSS WL0[136] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7285 VSS WL0[136] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7286 VSS WL0[136] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7287 VSS WL0[136] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7288 VSS WL0[136] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7289 VSS WL0[136] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7290 VSS WL0[136] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7291 VSS WL0[136] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7292 VSS WL0[136] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7293 VSS WL0[136] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7294 VSS WL0[136] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7295 VSS WL0[136] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7296 VSS WL0[136] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7297 VSS WL0[136] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7298 VSS WL0[136] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7299 VSS WL0[136] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7300 VSS WL0[136] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7301 VSS WL0[136] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7302 VSS WL0[136] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7303 VSS WL0[136] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7304 VSS WL0[136] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7305 VSS WL0[136] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7306 VSS WL0[136] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7307 VSS WL0[136] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7308 VSS WL0[136] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x890
XM7309 VSS WL0[137] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7310 VSS WL0[137] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7311 VSS WL0[137] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7312 VSS WL0[137] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7313 VSS WL0[137] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7314 VSS WL0[137] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7315 VSS WL0[137] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7316 VSS WL0[137] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7317 VSS WL0[137] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7318 VSS WL0[137] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7319 VSS WL0[137] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7320 VSS WL0[137] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7321 VSS WL0[137] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7322 VSS WL0[137] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7323 VSS WL0[137] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7324 VSS WL0[137] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7325 VSS WL0[137] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7326 VSS WL0[137] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7327 VSS WL0[137] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7328 VSS WL0[137] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7329 VSS WL0[137] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7330 VSS WL0[137] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7331 VSS WL0[137] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7332 VSS WL0[137] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7333 VSS WL0[137] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7334 VSS WL0[137] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7335 VSS WL0[137] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7336 VSS WL0[137] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7337 VSS WL0[137] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7338 VSS WL0[137] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7339 VSS WL0[137] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7340 VSS WL0[137] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7341 VSS WL0[137] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7342 VSS WL0[137] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7343 VSS WL0[137] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7344 VSS WL0[137] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7345 VSS WL0[137] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7346 VSS WL0[137] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7347 VSS WL0[137] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7348 VSS WL0[137] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7349 VSS WL0[137] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7350 VSS WL0[137] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7351 VSS WL0[137] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7352 VSS WL0[137] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7353 VSS WL0[137] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7354 VSS WL0[137] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7355 VSS WL0[137] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7356 VSS WL0[137] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7357 VSS WL0[137] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7358 VSS WL0[137] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7359 VSS WL0[137] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7360 VSS WL0[137] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7361 VSS WL0[137] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7362 VSS WL0[137] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7363 VSS WL0[137] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7364 VSS WL0[137] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7365 VSS WL0[137] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7366 VSS WL0[137] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7367 VSS WL0[137] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7368 VSS WL0[137] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7369 VSS WL0[137] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7370 VSS WL0[137] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7371 VSS WL0[137] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x8a0
XM7372 VSS WL0[138] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7373 VSS WL0[138] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7374 VSS WL0[138] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7375 VSS WL0[138] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7376 VSS WL0[138] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7377 VSS WL0[138] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7378 VSS WL0[138] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7379 VSS WL0[138] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7380 VSS WL0[138] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7381 VSS WL0[138] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7382 VSS WL0[138] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7383 VSS WL0[138] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7384 VSS WL0[138] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7385 VSS WL0[138] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7386 VSS WL0[138] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7387 VSS WL0[138] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7388 VSS WL0[138] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7389 VSS WL0[138] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7390 VSS WL0[138] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7391 VSS WL0[138] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7392 VSS WL0[138] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7393 VSS WL0[138] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7394 VSS WL0[138] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7395 VSS WL0[138] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7396 VSS WL0[138] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7397 VSS WL0[138] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7398 VSS WL0[138] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7399 VSS WL0[138] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7400 VSS WL0[138] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7401 VSS WL0[138] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7402 VSS WL0[138] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7403 VSS WL0[138] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7404 VSS WL0[138] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7405 VSS WL0[138] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7406 VSS WL0[138] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7407 VSS WL0[138] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7408 VSS WL0[138] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7409 VSS WL0[138] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7410 VSS WL0[138] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7411 VSS WL0[138] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7412 VSS WL0[138] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7413 VSS WL0[138] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7414 VSS WL0[138] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7415 VSS WL0[138] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7416 VSS WL0[138] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7417 VSS WL0[138] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7418 VSS WL0[138] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7419 VSS WL0[138] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7420 VSS WL0[138] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7421 VSS WL0[138] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7422 VSS WL0[138] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7423 VSS WL0[138] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x8b0
XM7424 VSS WL0[139] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7425 VSS WL0[139] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7426 VSS WL0[139] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7427 VSS WL0[139] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7428 VSS WL0[139] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7429 VSS WL0[139] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7430 VSS WL0[139] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7431 VSS WL0[139] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7432 VSS WL0[139] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7433 VSS WL0[139] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7434 VSS WL0[139] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7435 VSS WL0[139] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7436 VSS WL0[139] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7437 VSS WL0[139] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7438 VSS WL0[139] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7439 VSS WL0[139] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7440 VSS WL0[139] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7441 VSS WL0[139] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7442 VSS WL0[139] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7443 VSS WL0[139] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7444 VSS WL0[139] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7445 VSS WL0[139] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7446 VSS WL0[139] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7447 VSS WL0[139] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7448 VSS WL0[139] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7449 VSS WL0[139] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7450 VSS WL0[139] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7451 VSS WL0[139] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7452 VSS WL0[139] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7453 VSS WL0[139] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7454 VSS WL0[139] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7455 VSS WL0[139] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7456 VSS WL0[139] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7457 VSS WL0[139] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7458 VSS WL0[139] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7459 VSS WL0[139] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7460 VSS WL0[139] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7461 VSS WL0[139] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7462 VSS WL0[139] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7463 VSS WL0[139] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7464 VSS WL0[139] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7465 VSS WL0[139] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7466 VSS WL0[139] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7467 VSS WL0[139] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7468 VSS WL0[139] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7469 VSS WL0[139] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7470 VSS WL0[139] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7471 VSS WL0[139] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7472 VSS WL0[139] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7473 VSS WL0[139] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7474 VSS WL0[139] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7475 VSS WL0[139] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7476 VSS WL0[139] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7477 VSS WL0[139] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7478 VSS WL0[139] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7479 VSS WL0[139] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7480 VSS WL0[139] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7481 VSS WL0[139] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7482 VSS WL0[139] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7483 VSS WL0[139] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7484 VSS WL0[139] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7485 VSS WL0[139] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7486 VSS WL0[139] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7487 VSS WL0[139] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7488 VSS WL0[139] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7489 VSS WL0[139] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7490 VSS WL0[139] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7491 VSS WL0[139] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x8c0
XM7492 VSS WL0[140] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7493 VSS WL0[140] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7494 VSS WL0[140] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7495 VSS WL0[140] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7496 VSS WL0[140] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7497 VSS WL0[140] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7498 VSS WL0[140] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7499 VSS WL0[140] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7500 VSS WL0[140] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7501 VSS WL0[140] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7502 VSS WL0[140] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7503 VSS WL0[140] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7504 VSS WL0[140] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7505 VSS WL0[140] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7506 VSS WL0[140] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7507 VSS WL0[140] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7508 VSS WL0[140] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7509 VSS WL0[140] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7510 VSS WL0[140] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7511 VSS WL0[140] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7512 VSS WL0[140] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7513 VSS WL0[140] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7514 VSS WL0[140] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7515 VSS WL0[140] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7516 VSS WL0[140] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7517 VSS WL0[140] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7518 VSS WL0[140] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7519 VSS WL0[140] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7520 VSS WL0[140] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7521 VSS WL0[140] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7522 VSS WL0[140] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7523 VSS WL0[140] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7524 VSS WL0[140] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7525 VSS WL0[140] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7526 VSS WL0[140] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7527 VSS WL0[140] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7528 VSS WL0[140] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7529 VSS WL0[140] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7530 VSS WL0[140] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7531 VSS WL0[140] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7532 VSS WL0[140] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7533 VSS WL0[140] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7534 VSS WL0[140] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7535 VSS WL0[140] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7536 VSS WL0[140] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7537 VSS WL0[140] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7538 VSS WL0[140] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7539 VSS WL0[140] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7540 VSS WL0[140] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7541 VSS WL0[140] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7542 VSS WL0[140] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7543 VSS WL0[140] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7544 VSS WL0[140] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7545 VSS WL0[140] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7546 VSS WL0[140] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7547 VSS WL0[140] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7548 VSS WL0[140] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7549 VSS WL0[140] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7550 VSS WL0[140] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7551 VSS WL0[140] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7552 VSS WL0[140] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7553 VSS WL0[140] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x8d0
XM7554 VSS WL0[141] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7555 VSS WL0[141] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7556 VSS WL0[141] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7557 VSS WL0[141] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7558 VSS WL0[141] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7559 VSS WL0[141] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7560 VSS WL0[141] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7561 VSS WL0[141] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7562 VSS WL0[141] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7563 VSS WL0[141] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7564 VSS WL0[141] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7565 VSS WL0[141] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7566 VSS WL0[141] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7567 VSS WL0[141] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7568 VSS WL0[141] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7569 VSS WL0[141] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7570 VSS WL0[141] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7571 VSS WL0[141] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7572 VSS WL0[141] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7573 VSS WL0[141] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7574 VSS WL0[141] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7575 VSS WL0[141] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7576 VSS WL0[141] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7577 VSS WL0[141] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7578 VSS WL0[141] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7579 VSS WL0[141] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7580 VSS WL0[141] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7581 VSS WL0[141] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7582 VSS WL0[141] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7583 VSS WL0[141] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7584 VSS WL0[141] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7585 VSS WL0[141] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7586 VSS WL0[141] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7587 VSS WL0[141] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7588 VSS WL0[141] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7589 VSS WL0[141] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7590 VSS WL0[141] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7591 VSS WL0[141] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7592 VSS WL0[141] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7593 VSS WL0[141] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7594 VSS WL0[141] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7595 VSS WL0[141] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7596 VSS WL0[141] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7597 VSS WL0[141] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7598 VSS WL0[141] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7599 VSS WL0[141] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7600 VSS WL0[141] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7601 VSS WL0[141] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7602 VSS WL0[141] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7603 VSS WL0[141] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7604 VSS WL0[141] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x8e0
XM7605 VSS WL0[142] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7606 VSS WL0[142] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7607 VSS WL0[142] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7608 VSS WL0[142] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7609 VSS WL0[142] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7610 VSS WL0[142] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7611 VSS WL0[142] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7612 VSS WL0[142] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7613 VSS WL0[142] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7614 VSS WL0[142] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7615 VSS WL0[142] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7616 VSS WL0[142] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7617 VSS WL0[142] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7618 VSS WL0[142] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7619 VSS WL0[142] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7620 VSS WL0[142] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7621 VSS WL0[142] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7622 VSS WL0[142] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7623 VSS WL0[142] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7624 VSS WL0[142] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7625 VSS WL0[142] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7626 VSS WL0[142] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7627 VSS WL0[142] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7628 VSS WL0[142] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7629 VSS WL0[142] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7630 VSS WL0[142] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7631 VSS WL0[142] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7632 VSS WL0[142] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7633 VSS WL0[142] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7634 VSS WL0[142] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7635 VSS WL0[142] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7636 VSS WL0[142] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7637 VSS WL0[142] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7638 VSS WL0[142] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7639 VSS WL0[142] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7640 VSS WL0[142] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7641 VSS WL0[142] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7642 VSS WL0[142] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7643 VSS WL0[142] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7644 VSS WL0[142] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7645 VSS WL0[142] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7646 VSS WL0[142] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7647 VSS WL0[142] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7648 VSS WL0[142] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7649 VSS WL0[142] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7650 VSS WL0[142] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7651 VSS WL0[142] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7652 VSS WL0[142] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7653 VSS WL0[142] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x8f0
XM7654 VSS WL0[143] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7655 VSS WL0[143] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7656 VSS WL0[143] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7657 VSS WL0[143] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7658 VSS WL0[143] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7659 VSS WL0[143] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7660 VSS WL0[143] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7661 VSS WL0[143] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7662 VSS WL0[143] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7663 VSS WL0[143] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7664 VSS WL0[143] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7665 VSS WL0[143] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7666 VSS WL0[143] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7667 VSS WL0[143] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7668 VSS WL0[143] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7669 VSS WL0[143] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7670 VSS WL0[143] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7671 VSS WL0[143] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7672 VSS WL0[143] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7673 VSS WL0[143] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7674 VSS WL0[143] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7675 VSS WL0[143] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7676 VSS WL0[143] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7677 VSS WL0[143] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7678 VSS WL0[143] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7679 VSS WL0[143] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7680 VSS WL0[143] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7681 VSS WL0[143] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7682 VSS WL0[143] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7683 VSS WL0[143] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7684 VSS WL0[143] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7685 VSS WL0[143] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7686 VSS WL0[143] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7687 VSS WL0[143] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7688 VSS WL0[143] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7689 VSS WL0[143] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7690 VSS WL0[143] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7691 VSS WL0[143] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7692 VSS WL0[143] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7693 VSS WL0[143] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7694 VSS WL0[143] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7695 VSS WL0[143] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7696 VSS WL0[143] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7697 VSS WL0[143] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7698 VSS WL0[143] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7699 VSS WL0[143] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7700 VSS WL0[143] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7701 VSS WL0[143] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7702 VSS WL0[143] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7703 VSS WL0[143] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7704 VSS WL0[143] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7705 VSS WL0[143] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7706 VSS WL0[143] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7707 VSS WL0[143] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7708 VSS WL0[143] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x900
XM7709 VSS WL0[144] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7710 VSS WL0[144] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7711 VSS WL0[144] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7712 VSS WL0[144] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7713 VSS WL0[144] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7714 VSS WL0[144] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7715 VSS WL0[144] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7716 VSS WL0[144] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7717 VSS WL0[144] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7718 VSS WL0[144] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7719 VSS WL0[144] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7720 VSS WL0[144] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7721 VSS WL0[144] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7722 VSS WL0[144] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7723 VSS WL0[144] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7724 VSS WL0[144] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7725 VSS WL0[144] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7726 VSS WL0[144] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7727 VSS WL0[144] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7728 VSS WL0[144] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7729 VSS WL0[144] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7730 VSS WL0[144] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7731 VSS WL0[144] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7732 VSS WL0[144] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7733 VSS WL0[144] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7734 VSS WL0[144] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7735 VSS WL0[144] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7736 VSS WL0[144] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7737 VSS WL0[144] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7738 VSS WL0[144] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7739 VSS WL0[144] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7740 VSS WL0[144] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7741 VSS WL0[144] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7742 VSS WL0[144] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7743 VSS WL0[144] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7744 VSS WL0[144] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7745 VSS WL0[144] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7746 VSS WL0[144] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7747 VSS WL0[144] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7748 VSS WL0[144] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7749 VSS WL0[144] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7750 VSS WL0[144] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7751 VSS WL0[144] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7752 VSS WL0[144] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7753 VSS WL0[144] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7754 VSS WL0[144] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7755 VSS WL0[144] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7756 VSS WL0[144] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7757 VSS WL0[144] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7758 VSS WL0[144] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7759 VSS WL0[144] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7760 VSS WL0[144] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x910
XM7761 VSS WL0[145] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7762 VSS WL0[145] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7763 VSS WL0[145] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7764 VSS WL0[145] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7765 VSS WL0[145] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7766 VSS WL0[145] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7767 VSS WL0[145] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7768 VSS WL0[145] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7769 VSS WL0[145] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7770 VSS WL0[145] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7771 VSS WL0[145] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7772 VSS WL0[145] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7773 VSS WL0[145] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7774 VSS WL0[145] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7775 VSS WL0[145] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7776 VSS WL0[145] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7777 VSS WL0[145] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7778 VSS WL0[145] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7779 VSS WL0[145] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7780 VSS WL0[145] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7781 VSS WL0[145] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7782 VSS WL0[145] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7783 VSS WL0[145] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7784 VSS WL0[145] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7785 VSS WL0[145] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7786 VSS WL0[145] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7787 VSS WL0[145] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7788 VSS WL0[145] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7789 VSS WL0[145] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7790 VSS WL0[145] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7791 VSS WL0[145] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7792 VSS WL0[145] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7793 VSS WL0[145] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7794 VSS WL0[145] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7795 VSS WL0[145] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7796 VSS WL0[145] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7797 VSS WL0[145] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7798 VSS WL0[145] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7799 VSS WL0[145] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7800 VSS WL0[145] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7801 VSS WL0[145] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7802 VSS WL0[145] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7803 VSS WL0[145] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7804 VSS WL0[145] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7805 VSS WL0[145] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7806 VSS WL0[145] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7807 VSS WL0[145] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7808 VSS WL0[145] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7809 VSS WL0[145] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7810 VSS WL0[145] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7811 VSS WL0[145] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7812 VSS WL0[145] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x920
XM7813 VSS WL0[146] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7814 VSS WL0[146] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7815 VSS WL0[146] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7816 VSS WL0[146] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7817 VSS WL0[146] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7818 VSS WL0[146] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7819 VSS WL0[146] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7820 VSS WL0[146] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7821 VSS WL0[146] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7822 VSS WL0[146] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7823 VSS WL0[146] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7824 VSS WL0[146] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7825 VSS WL0[146] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7826 VSS WL0[146] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7827 VSS WL0[146] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7828 VSS WL0[146] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7829 VSS WL0[146] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7830 VSS WL0[146] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7831 VSS WL0[146] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7832 VSS WL0[146] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7833 VSS WL0[146] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7834 VSS WL0[146] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7835 VSS WL0[146] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7836 VSS WL0[146] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7837 VSS WL0[146] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7838 VSS WL0[146] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7839 VSS WL0[146] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7840 VSS WL0[146] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7841 VSS WL0[146] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7842 VSS WL0[146] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7843 VSS WL0[146] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7844 VSS WL0[146] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7845 VSS WL0[146] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7846 VSS WL0[146] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7847 VSS WL0[146] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7848 VSS WL0[146] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7849 VSS WL0[146] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7850 VSS WL0[146] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7851 VSS WL0[146] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7852 VSS WL0[146] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7853 VSS WL0[146] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7854 VSS WL0[146] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7855 VSS WL0[146] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7856 VSS WL0[146] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7857 VSS WL0[146] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7858 VSS WL0[146] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7859 VSS WL0[146] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7860 VSS WL0[146] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7861 VSS WL0[146] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7862 VSS WL0[146] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7863 VSS WL0[146] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7864 VSS WL0[146] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7865 VSS WL0[146] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7866 VSS WL0[146] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x930
XM7867 VSS WL0[147] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7868 VSS WL0[147] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7869 VSS WL0[147] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7870 VSS WL0[147] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7871 VSS WL0[147] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7872 VSS WL0[147] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7873 VSS WL0[147] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7874 VSS WL0[147] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7875 VSS WL0[147] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7876 VSS WL0[147] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7877 VSS WL0[147] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7878 VSS WL0[147] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7879 VSS WL0[147] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7880 VSS WL0[147] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7881 VSS WL0[147] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7882 VSS WL0[147] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7883 VSS WL0[147] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7884 VSS WL0[147] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7885 VSS WL0[147] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7886 VSS WL0[147] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7887 VSS WL0[147] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7888 VSS WL0[147] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7889 VSS WL0[147] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7890 VSS WL0[147] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7891 VSS WL0[147] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7892 VSS WL0[147] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7893 VSS WL0[147] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7894 VSS WL0[147] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7895 VSS WL0[147] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7896 VSS WL0[147] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7897 VSS WL0[147] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7898 VSS WL0[147] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7899 VSS WL0[147] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7900 VSS WL0[147] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7901 VSS WL0[147] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7902 VSS WL0[147] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7903 VSS WL0[147] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7904 VSS WL0[147] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7905 VSS WL0[147] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7906 VSS WL0[147] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7907 VSS WL0[147] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7908 VSS WL0[147] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7909 VSS WL0[147] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7910 VSS WL0[147] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7911 VSS WL0[147] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7912 VSS WL0[147] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7913 VSS WL0[147] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7914 VSS WL0[147] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7915 VSS WL0[147] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7916 VSS WL0[147] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7917 VSS WL0[147] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7918 VSS WL0[147] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7919 VSS WL0[147] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x940
XM7920 VSS WL0[148] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7921 VSS WL0[148] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7922 VSS WL0[148] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7923 VSS WL0[148] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7924 VSS WL0[148] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7925 VSS WL0[148] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7926 VSS WL0[148] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7927 VSS WL0[148] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7928 VSS WL0[148] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7929 VSS WL0[148] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7930 VSS WL0[148] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7931 VSS WL0[148] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7932 VSS WL0[148] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7933 VSS WL0[148] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7934 VSS WL0[148] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7935 VSS WL0[148] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7936 VSS WL0[148] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7937 VSS WL0[148] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7938 VSS WL0[148] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7939 VSS WL0[148] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7940 VSS WL0[148] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7941 VSS WL0[148] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7942 VSS WL0[148] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7943 VSS WL0[148] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7944 VSS WL0[148] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7945 VSS WL0[148] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7946 VSS WL0[148] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7947 VSS WL0[148] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7948 VSS WL0[148] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7949 VSS WL0[148] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7950 VSS WL0[148] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7951 VSS WL0[148] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7952 VSS WL0[148] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7953 VSS WL0[148] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7954 VSS WL0[148] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7955 VSS WL0[148] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7956 VSS WL0[148] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7957 VSS WL0[148] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7958 VSS WL0[148] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7959 VSS WL0[148] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7960 VSS WL0[148] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7961 VSS WL0[148] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7962 VSS WL0[148] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7963 VSS WL0[148] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7964 VSS WL0[148] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x950
XM7965 VSS WL0[149] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7966 VSS WL0[149] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7967 VSS WL0[149] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7968 VSS WL0[149] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7969 VSS WL0[149] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7970 VSS WL0[149] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7971 VSS WL0[149] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7972 VSS WL0[149] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7973 VSS WL0[149] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7974 VSS WL0[149] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7975 VSS WL0[149] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7976 VSS WL0[149] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7977 VSS WL0[149] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7978 VSS WL0[149] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7979 VSS WL0[149] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7980 VSS WL0[149] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7981 VSS WL0[149] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7982 VSS WL0[149] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7983 VSS WL0[149] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7984 VSS WL0[149] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7985 VSS WL0[149] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7986 VSS WL0[149] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7987 VSS WL0[149] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7988 VSS WL0[149] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7989 VSS WL0[149] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7990 VSS WL0[149] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7991 VSS WL0[149] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7992 VSS WL0[149] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7993 VSS WL0[149] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7994 VSS WL0[149] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7995 VSS WL0[149] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7996 VSS WL0[149] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7997 VSS WL0[149] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7998 VSS WL0[149] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM7999 VSS WL0[149] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8000 VSS WL0[149] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8001 VSS WL0[149] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8002 VSS WL0[149] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8003 VSS WL0[149] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8004 VSS WL0[149] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x960
XM8005 VSS WL0[150] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8006 VSS WL0[150] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8007 VSS WL0[150] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8008 VSS WL0[150] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8009 VSS WL0[150] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8010 VSS WL0[150] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8011 VSS WL0[150] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8012 VSS WL0[150] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8013 VSS WL0[150] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8014 VSS WL0[150] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8015 VSS WL0[150] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8016 VSS WL0[150] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8017 VSS WL0[150] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8018 VSS WL0[150] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8019 VSS WL0[150] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8020 VSS WL0[150] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x970
XM8021 VSS WL0[151] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8022 VSS WL0[151] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8023 VSS WL0[151] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8024 VSS WL0[151] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8025 VSS WL0[151] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8026 VSS WL0[151] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8027 VSS WL0[151] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8028 VSS WL0[151] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8029 VSS WL0[151] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8030 VSS WL0[151] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8031 VSS WL0[151] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8032 VSS WL0[151] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8033 VSS WL0[151] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8034 VSS WL0[151] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8035 VSS WL0[151] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8036 VSS WL0[151] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8037 VSS WL0[151] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8038 VSS WL0[151] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8039 VSS WL0[151] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8040 VSS WL0[151] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x980
XM8041 VSS WL0[152] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8042 VSS WL0[152] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8043 VSS WL0[152] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8044 VSS WL0[152] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8045 VSS WL0[152] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8046 VSS WL0[152] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8047 VSS WL0[152] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8048 VSS WL0[152] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8049 VSS WL0[152] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8050 VSS WL0[152] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8051 VSS WL0[152] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8052 VSS WL0[152] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8053 VSS WL0[152] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8054 VSS WL0[152] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8055 VSS WL0[152] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8056 VSS WL0[152] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8057 VSS WL0[152] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8058 VSS WL0[152] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8059 VSS WL0[152] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8060 VSS WL0[152] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x990
XM8061 VSS WL0[153] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8062 VSS WL0[153] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8063 VSS WL0[153] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8064 VSS WL0[153] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8065 VSS WL0[153] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8066 VSS WL0[153] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8067 VSS WL0[153] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8068 VSS WL0[153] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8069 VSS WL0[153] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8070 VSS WL0[153] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8071 VSS WL0[153] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8072 VSS WL0[153] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8073 VSS WL0[153] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8074 VSS WL0[153] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8075 VSS WL0[153] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8076 VSS WL0[153] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8077 VSS WL0[153] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8078 VSS WL0[153] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8079 VSS WL0[153] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x9a0
XM8080 VSS WL0[154] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8081 VSS WL0[154] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8082 VSS WL0[154] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8083 VSS WL0[154] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8084 VSS WL0[154] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8085 VSS WL0[154] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8086 VSS WL0[154] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8087 VSS WL0[154] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8088 VSS WL0[154] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8089 VSS WL0[154] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8090 VSS WL0[154] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8091 VSS WL0[154] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8092 VSS WL0[154] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8093 VSS WL0[154] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8094 VSS WL0[154] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8095 VSS WL0[154] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8096 VSS WL0[154] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8097 VSS WL0[154] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8098 VSS WL0[154] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8099 VSS WL0[154] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x9b0
XM8100 VSS WL0[155] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8101 VSS WL0[155] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8102 VSS WL0[155] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8103 VSS WL0[155] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8104 VSS WL0[155] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8105 VSS WL0[155] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8106 VSS WL0[155] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8107 VSS WL0[155] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8108 VSS WL0[155] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8109 VSS WL0[155] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8110 VSS WL0[155] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8111 VSS WL0[155] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8112 VSS WL0[155] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8113 VSS WL0[155] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8114 VSS WL0[155] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8115 VSS WL0[155] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8116 VSS WL0[155] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8117 VSS WL0[155] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x9c0
XM8118 VSS WL0[156] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8119 VSS WL0[156] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8120 VSS WL0[156] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8121 VSS WL0[156] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8122 VSS WL0[156] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8123 VSS WL0[156] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8124 VSS WL0[156] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8125 VSS WL0[156] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8126 VSS WL0[156] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8127 VSS WL0[156] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8128 VSS WL0[156] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8129 VSS WL0[156] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8130 VSS WL0[156] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8131 VSS WL0[156] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8132 VSS WL0[156] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8133 VSS WL0[156] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8134 VSS WL0[156] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8135 VSS WL0[156] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8136 VSS WL0[156] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8137 VSS WL0[156] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8138 VSS WL0[156] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8139 VSS WL0[156] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8140 VSS WL0[156] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8141 VSS WL0[156] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x9d0
XM8142 VSS WL0[157] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8143 VSS WL0[157] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8144 VSS WL0[157] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8145 VSS WL0[157] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8146 VSS WL0[157] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8147 VSS WL0[157] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8148 VSS WL0[157] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8149 VSS WL0[157] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8150 VSS WL0[157] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8151 VSS WL0[157] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8152 VSS WL0[157] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8153 VSS WL0[157] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8154 VSS WL0[157] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8155 VSS WL0[157] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8156 VSS WL0[157] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8157 VSS WL0[157] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8158 VSS WL0[157] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8159 VSS WL0[157] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8160 VSS WL0[157] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8161 VSS WL0[157] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8162 VSS WL0[157] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8163 VSS WL0[157] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8164 VSS WL0[157] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8165 VSS WL0[157] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x9e0
XM8166 VSS WL0[158] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8167 VSS WL0[158] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8168 VSS WL0[158] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8169 VSS WL0[158] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8170 VSS WL0[158] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8171 VSS WL0[158] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8172 VSS WL0[158] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8173 VSS WL0[158] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8174 VSS WL0[158] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8175 VSS WL0[158] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8176 VSS WL0[158] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8177 VSS WL0[158] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8178 VSS WL0[158] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8179 VSS WL0[158] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8180 VSS WL0[158] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8181 VSS WL0[158] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8182 VSS WL0[158] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8183 VSS WL0[158] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8184 VSS WL0[158] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8185 VSS WL0[158] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8186 VSS WL0[158] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8187 VSS WL0[158] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8188 VSS WL0[158] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8189 VSS WL0[158] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0x9f0
XM8190 VSS WL0[159] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8191 VSS WL0[159] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8192 VSS WL0[159] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8193 VSS WL0[159] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8194 VSS WL0[159] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8195 VSS WL0[159] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8196 VSS WL0[159] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8197 VSS WL0[159] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8198 VSS WL0[159] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8199 VSS WL0[159] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8200 VSS WL0[159] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8201 VSS WL0[159] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8202 VSS WL0[159] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8203 VSS WL0[159] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8204 VSS WL0[159] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8205 VSS WL0[159] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8206 VSS WL0[159] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8207 VSS WL0[159] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8208 VSS WL0[159] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8209 VSS WL0[159] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8210 VSS WL0[159] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8211 VSS WL0[159] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* addr: 0xa00
XM8212 VSS WL0[160] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8213 VSS WL0[160] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8214 VSS WL0[160] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8215 VSS WL0[160] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8216 VSS WL0[160] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8217 VSS WL0[160] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8218 VSS WL0[160] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8219 VSS WL0[160] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8220 VSS WL0[160] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8221 VSS WL0[160] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8222 VSS WL0[160] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8223 VSS WL0[160] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8224 VSS WL0[160] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8225 VSS WL0[160] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8226 VSS WL0[160] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8227 VSS WL0[160] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8228 VSS WL0[160] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8229 VSS WL0[160] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8230 VSS WL0[160] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8231 VSS WL0[160] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8232 VSS WL0[160] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8233 VSS WL0[160] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8234 VSS WL0[160] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8235 VSS WL0[160] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8236 VSS WL0[160] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XM8237 VSS WL0[160] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
* Read muxers
XRDn[0] RD_M[0] COL_B10_p[0] BL[0] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[0] RD_M[0] COL_B10_n[0] BL[0] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[1] RD_M[1] COL_B10_p[0] BL[1] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[1] RD_M[1] COL_B10_n[0] BL[1] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[2] RD_M[2] COL_B10_p[0] BL[2] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[2] RD_M[2] COL_B10_n[0] BL[2] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[3] RD_M[3] COL_B10_p[0] BL[3] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[3] RD_M[3] COL_B10_n[0] BL[3] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[4] RD_M[4] COL_B10_p[0] BL[4] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[4] RD_M[4] COL_B10_n[0] BL[4] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[5] RD_M[5] COL_B10_p[0] BL[5] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[5] RD_M[5] COL_B10_n[0] BL[5] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[6] RD_M[6] COL_B10_p[0] BL[6] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[6] RD_M[6] COL_B10_n[0] BL[6] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[7] RD_M[7] COL_B10_p[0] BL[7] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[7] RD_M[7] COL_B10_n[0] BL[7] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[8] RD_M[8] COL_B11_p[0] BL[8] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[8] RD_M[8] COL_B11_n[0] BL[8] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[9] RD_M[9] COL_B11_p[0] BL[9] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[9] RD_M[9] COL_B11_n[0] BL[9] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[10] RD_M[10] COL_B11_p[0] BL[10] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[10] RD_M[10] COL_B11_n[0] BL[10] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[11] RD_M[11] COL_B11_p[0] BL[11] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[11] RD_M[11] COL_B11_n[0] BL[11] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[12] RD_M[12] COL_B11_p[0] BL[12] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[12] RD_M[12] COL_B11_n[0] BL[12] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[13] RD_M[13] COL_B11_p[0] BL[13] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[13] RD_M[13] COL_B11_n[0] BL[13] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[14] RD_M[14] COL_B11_p[0] BL[14] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[14] RD_M[14] COL_B11_n[0] BL[14] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[15] RD_M[15] COL_B11_p[0] BL[15] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[15] RD_M[15] COL_B11_n[0] BL[15] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[16] RD_M[16] COL_B12_p[0] BL[16] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[16] RD_M[16] COL_B12_n[0] BL[16] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[17] RD_M[17] COL_B12_p[0] BL[17] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[17] RD_M[17] COL_B12_n[0] BL[17] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[18] RD_M[18] COL_B12_p[0] BL[18] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[18] RD_M[18] COL_B12_n[0] BL[18] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[19] RD_M[19] COL_B12_p[0] BL[19] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[19] RD_M[19] COL_B12_n[0] BL[19] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[20] RD_M[20] COL_B12_p[0] BL[20] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[20] RD_M[20] COL_B12_n[0] BL[20] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[21] RD_M[21] COL_B12_p[0] BL[21] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[21] RD_M[21] COL_B12_n[0] BL[21] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[22] RD_M[22] COL_B12_p[0] BL[22] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[22] RD_M[22] COL_B12_n[0] BL[22] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[23] RD_M[23] COL_B12_p[0] BL[23] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[23] RD_M[23] COL_B12_n[0] BL[23] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[24] RD_M[24] COL_B13_p[0] BL[24] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[24] RD_M[24] COL_B13_n[0] BL[24] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[25] RD_M[25] COL_B13_p[0] BL[25] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[25] RD_M[25] COL_B13_n[0] BL[25] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[26] RD_M[26] COL_B13_p[0] BL[26] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[26] RD_M[26] COL_B13_n[0] BL[26] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[27] RD_M[27] COL_B13_p[0] BL[27] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[27] RD_M[27] COL_B13_n[0] BL[27] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[28] RD_M[28] COL_B13_p[0] BL[28] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[28] RD_M[28] COL_B13_n[0] BL[28] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[29] RD_M[29] COL_B13_p[0] BL[29] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[29] RD_M[29] COL_B13_n[0] BL[29] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[30] RD_M[30] COL_B13_p[0] BL[30] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[30] RD_M[30] COL_B13_n[0] BL[30] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[31] RD_M[31] COL_B13_p[0] BL[31] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[31] RD_M[31] COL_B13_n[0] BL[31] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[32] RD_M[0] COL_B10_p[1] BL[32] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[32] RD_M[0] COL_B10_n[1] BL[32] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[33] RD_M[1] COL_B10_p[1] BL[33] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[33] RD_M[1] COL_B10_n[1] BL[33] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[34] RD_M[2] COL_B10_p[1] BL[34] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[34] RD_M[2] COL_B10_n[1] BL[34] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[35] RD_M[3] COL_B10_p[1] BL[35] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[35] RD_M[3] COL_B10_n[1] BL[35] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[36] RD_M[4] COL_B10_p[1] BL[36] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[36] RD_M[4] COL_B10_n[1] BL[36] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[37] RD_M[5] COL_B10_p[1] BL[37] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[37] RD_M[5] COL_B10_n[1] BL[37] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[38] RD_M[6] COL_B10_p[1] BL[38] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[38] RD_M[6] COL_B10_n[1] BL[38] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[39] RD_M[7] COL_B10_p[1] BL[39] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[39] RD_M[7] COL_B10_n[1] BL[39] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[40] RD_M[8] COL_B11_p[1] BL[40] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[40] RD_M[8] COL_B11_n[1] BL[40] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[41] RD_M[9] COL_B11_p[1] BL[41] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[41] RD_M[9] COL_B11_n[1] BL[41] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[42] RD_M[10] COL_B11_p[1] BL[42] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[42] RD_M[10] COL_B11_n[1] BL[42] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[43] RD_M[11] COL_B11_p[1] BL[43] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[43] RD_M[11] COL_B11_n[1] BL[43] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[44] RD_M[12] COL_B11_p[1] BL[44] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[44] RD_M[12] COL_B11_n[1] BL[44] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[45] RD_M[13] COL_B11_p[1] BL[45] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[45] RD_M[13] COL_B11_n[1] BL[45] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[46] RD_M[14] COL_B11_p[1] BL[46] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[46] RD_M[14] COL_B11_n[1] BL[46] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[47] RD_M[15] COL_B11_p[1] BL[47] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[47] RD_M[15] COL_B11_n[1] BL[47] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[48] RD_M[16] COL_B12_p[1] BL[48] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[48] RD_M[16] COL_B12_n[1] BL[48] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[49] RD_M[17] COL_B12_p[1] BL[49] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[49] RD_M[17] COL_B12_n[1] BL[49] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[50] RD_M[18] COL_B12_p[1] BL[50] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[50] RD_M[18] COL_B12_n[1] BL[50] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[51] RD_M[19] COL_B12_p[1] BL[51] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[51] RD_M[19] COL_B12_n[1] BL[51] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[52] RD_M[20] COL_B12_p[1] BL[52] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[52] RD_M[20] COL_B12_n[1] BL[52] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[53] RD_M[21] COL_B12_p[1] BL[53] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[53] RD_M[21] COL_B12_n[1] BL[53] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[54] RD_M[22] COL_B12_p[1] BL[54] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[54] RD_M[22] COL_B12_n[1] BL[54] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[55] RD_M[23] COL_B12_p[1] BL[55] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[55] RD_M[23] COL_B12_n[1] BL[55] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[56] RD_M[24] COL_B13_p[1] BL[56] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[56] RD_M[24] COL_B13_n[1] BL[56] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[57] RD_M[25] COL_B13_p[1] BL[57] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[57] RD_M[25] COL_B13_n[1] BL[57] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[58] RD_M[26] COL_B13_p[1] BL[58] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[58] RD_M[26] COL_B13_n[1] BL[58] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[59] RD_M[27] COL_B13_p[1] BL[59] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[59] RD_M[27] COL_B13_n[1] BL[59] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[60] RD_M[28] COL_B13_p[1] BL[60] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[60] RD_M[28] COL_B13_n[1] BL[60] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[61] RD_M[29] COL_B13_p[1] BL[61] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[61] RD_M[29] COL_B13_n[1] BL[61] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[62] RD_M[30] COL_B13_p[1] BL[62] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[62] RD_M[30] COL_B13_n[1] BL[62] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[63] RD_M[31] COL_B13_p[1] BL[63] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[63] RD_M[31] COL_B13_n[1] BL[63] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[64] RD_M[0] COL_B10_p[2] BL[64] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[64] RD_M[0] COL_B10_n[2] BL[64] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[65] RD_M[1] COL_B10_p[2] BL[65] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[65] RD_M[1] COL_B10_n[2] BL[65] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[66] RD_M[2] COL_B10_p[2] BL[66] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[66] RD_M[2] COL_B10_n[2] BL[66] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[67] RD_M[3] COL_B10_p[2] BL[67] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[67] RD_M[3] COL_B10_n[2] BL[67] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[68] RD_M[4] COL_B10_p[2] BL[68] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[68] RD_M[4] COL_B10_n[2] BL[68] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[69] RD_M[5] COL_B10_p[2] BL[69] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[69] RD_M[5] COL_B10_n[2] BL[69] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[70] RD_M[6] COL_B10_p[2] BL[70] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[70] RD_M[6] COL_B10_n[2] BL[70] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[71] RD_M[7] COL_B10_p[2] BL[71] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[71] RD_M[7] COL_B10_n[2] BL[71] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[72] RD_M[8] COL_B11_p[2] BL[72] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[72] RD_M[8] COL_B11_n[2] BL[72] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[73] RD_M[9] COL_B11_p[2] BL[73] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[73] RD_M[9] COL_B11_n[2] BL[73] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[74] RD_M[10] COL_B11_p[2] BL[74] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[74] RD_M[10] COL_B11_n[2] BL[74] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[75] RD_M[11] COL_B11_p[2] BL[75] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[75] RD_M[11] COL_B11_n[2] BL[75] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[76] RD_M[12] COL_B11_p[2] BL[76] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[76] RD_M[12] COL_B11_n[2] BL[76] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[77] RD_M[13] COL_B11_p[2] BL[77] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[77] RD_M[13] COL_B11_n[2] BL[77] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[78] RD_M[14] COL_B11_p[2] BL[78] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[78] RD_M[14] COL_B11_n[2] BL[78] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[79] RD_M[15] COL_B11_p[2] BL[79] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[79] RD_M[15] COL_B11_n[2] BL[79] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[80] RD_M[16] COL_B12_p[2] BL[80] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[80] RD_M[16] COL_B12_n[2] BL[80] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[81] RD_M[17] COL_B12_p[2] BL[81] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[81] RD_M[17] COL_B12_n[2] BL[81] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[82] RD_M[18] COL_B12_p[2] BL[82] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[82] RD_M[18] COL_B12_n[2] BL[82] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[83] RD_M[19] COL_B12_p[2] BL[83] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[83] RD_M[19] COL_B12_n[2] BL[83] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[84] RD_M[20] COL_B12_p[2] BL[84] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[84] RD_M[20] COL_B12_n[2] BL[84] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[85] RD_M[21] COL_B12_p[2] BL[85] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[85] RD_M[21] COL_B12_n[2] BL[85] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[86] RD_M[22] COL_B12_p[2] BL[86] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[86] RD_M[22] COL_B12_n[2] BL[86] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[87] RD_M[23] COL_B12_p[2] BL[87] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[87] RD_M[23] COL_B12_n[2] BL[87] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[88] RD_M[24] COL_B13_p[2] BL[88] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[88] RD_M[24] COL_B13_n[2] BL[88] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[89] RD_M[25] COL_B13_p[2] BL[89] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[89] RD_M[25] COL_B13_n[2] BL[89] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[90] RD_M[26] COL_B13_p[2] BL[90] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[90] RD_M[26] COL_B13_n[2] BL[90] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[91] RD_M[27] COL_B13_p[2] BL[91] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[91] RD_M[27] COL_B13_n[2] BL[91] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[92] RD_M[28] COL_B13_p[2] BL[92] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[92] RD_M[28] COL_B13_n[2] BL[92] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[93] RD_M[29] COL_B13_p[2] BL[93] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[93] RD_M[29] COL_B13_n[2] BL[93] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[94] RD_M[30] COL_B13_p[2] BL[94] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[94] RD_M[30] COL_B13_n[2] BL[94] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[95] RD_M[31] COL_B13_p[2] BL[95] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[95] RD_M[31] COL_B13_n[2] BL[95] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[96] RD_M[0] COL_B10_p[3] BL[96] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[96] RD_M[0] COL_B10_n[3] BL[96] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[97] RD_M[1] COL_B10_p[3] BL[97] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[97] RD_M[1] COL_B10_n[3] BL[97] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[98] RD_M[2] COL_B10_p[3] BL[98] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[98] RD_M[2] COL_B10_n[3] BL[98] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[99] RD_M[3] COL_B10_p[3] BL[99] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[99] RD_M[3] COL_B10_n[3] BL[99] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[100] RD_M[4] COL_B10_p[3] BL[100] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[100] RD_M[4] COL_B10_n[3] BL[100] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[101] RD_M[5] COL_B10_p[3] BL[101] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[101] RD_M[5] COL_B10_n[3] BL[101] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[102] RD_M[6] COL_B10_p[3] BL[102] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[102] RD_M[6] COL_B10_n[3] BL[102] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[103] RD_M[7] COL_B10_p[3] BL[103] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[103] RD_M[7] COL_B10_n[3] BL[103] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[104] RD_M[8] COL_B11_p[3] BL[104] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[104] RD_M[8] COL_B11_n[3] BL[104] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[105] RD_M[9] COL_B11_p[3] BL[105] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[105] RD_M[9] COL_B11_n[3] BL[105] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[106] RD_M[10] COL_B11_p[3] BL[106] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[106] RD_M[10] COL_B11_n[3] BL[106] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[107] RD_M[11] COL_B11_p[3] BL[107] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[107] RD_M[11] COL_B11_n[3] BL[107] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[108] RD_M[12] COL_B11_p[3] BL[108] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[108] RD_M[12] COL_B11_n[3] BL[108] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[109] RD_M[13] COL_B11_p[3] BL[109] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[109] RD_M[13] COL_B11_n[3] BL[109] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[110] RD_M[14] COL_B11_p[3] BL[110] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[110] RD_M[14] COL_B11_n[3] BL[110] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[111] RD_M[15] COL_B11_p[3] BL[111] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[111] RD_M[15] COL_B11_n[3] BL[111] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[112] RD_M[16] COL_B12_p[3] BL[112] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[112] RD_M[16] COL_B12_n[3] BL[112] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[113] RD_M[17] COL_B12_p[3] BL[113] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[113] RD_M[17] COL_B12_n[3] BL[113] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[114] RD_M[18] COL_B12_p[3] BL[114] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[114] RD_M[18] COL_B12_n[3] BL[114] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[115] RD_M[19] COL_B12_p[3] BL[115] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[115] RD_M[19] COL_B12_n[3] BL[115] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[116] RD_M[20] COL_B12_p[3] BL[116] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[116] RD_M[20] COL_B12_n[3] BL[116] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[117] RD_M[21] COL_B12_p[3] BL[117] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[117] RD_M[21] COL_B12_n[3] BL[117] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[118] RD_M[22] COL_B12_p[3] BL[118] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[118] RD_M[22] COL_B12_n[3] BL[118] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[119] RD_M[23] COL_B12_p[3] BL[119] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[119] RD_M[23] COL_B12_n[3] BL[119] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[120] RD_M[24] COL_B13_p[3] BL[120] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[120] RD_M[24] COL_B13_n[3] BL[120] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[121] RD_M[25] COL_B13_p[3] BL[121] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[121] RD_M[25] COL_B13_n[3] BL[121] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[122] RD_M[26] COL_B13_p[3] BL[122] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[122] RD_M[26] COL_B13_n[3] BL[122] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[123] RD_M[27] COL_B13_p[3] BL[123] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[123] RD_M[27] COL_B13_n[3] BL[123] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[124] RD_M[28] COL_B13_p[3] BL[124] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[124] RD_M[28] COL_B13_n[3] BL[124] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[125] RD_M[29] COL_B13_p[3] BL[125] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[125] RD_M[29] COL_B13_n[3] BL[125] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[126] RD_M[30] COL_B13_p[3] BL[126] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[126] RD_M[30] COL_B13_n[3] BL[126] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
XRDn[127] RD_M[31] COL_B13_p[3] BL[127] VSS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
XRDp[127] RD_M[31] COL_B13_n[3] BL[127] VCC sky130_fd_pr__pfet_01v8_hvt w=1000000u l=150000u
* Out invertors
xRBUF[0] RD_M[0] VSS VSS VCC VCC RD[0] sky130_fd_sc_hd__inv_1
xRBUF[1] RD_M[1] VSS VSS VCC VCC RD[1] sky130_fd_sc_hd__inv_1
xRBUF[2] RD_M[2] VSS VSS VCC VCC RD[2] sky130_fd_sc_hd__inv_1
xRBUF[3] RD_M[3] VSS VSS VCC VCC RD[3] sky130_fd_sc_hd__inv_1
xRBUF[4] RD_M[4] VSS VSS VCC VCC RD[4] sky130_fd_sc_hd__inv_1
xRBUF[5] RD_M[5] VSS VSS VCC VCC RD[5] sky130_fd_sc_hd__inv_1
xRBUF[6] RD_M[6] VSS VSS VCC VCC RD[6] sky130_fd_sc_hd__inv_1
xRBUF[7] RD_M[7] VSS VSS VCC VCC RD[7] sky130_fd_sc_hd__inv_1
xRBUF[8] RD_M[8] VSS VSS VCC VCC RD[8] sky130_fd_sc_hd__inv_1
xRBUF[9] RD_M[9] VSS VSS VCC VCC RD[9] sky130_fd_sc_hd__inv_1
xRBUF[10] RD_M[10] VSS VSS VCC VCC RD[10] sky130_fd_sc_hd__inv_1
xRBUF[11] RD_M[11] VSS VSS VCC VCC RD[11] sky130_fd_sc_hd__inv_1
xRBUF[12] RD_M[12] VSS VSS VCC VCC RD[12] sky130_fd_sc_hd__inv_1
xRBUF[13] RD_M[13] VSS VSS VCC VCC RD[13] sky130_fd_sc_hd__inv_1
xRBUF[14] RD_M[14] VSS VSS VCC VCC RD[14] sky130_fd_sc_hd__inv_1
xRBUF[15] RD_M[15] VSS VSS VCC VCC RD[15] sky130_fd_sc_hd__inv_1
xRBUF[16] RD_M[16] VSS VSS VCC VCC RD[16] sky130_fd_sc_hd__inv_1
xRBUF[17] RD_M[17] VSS VSS VCC VCC RD[17] sky130_fd_sc_hd__inv_1
xRBUF[18] RD_M[18] VSS VSS VCC VCC RD[18] sky130_fd_sc_hd__inv_1
xRBUF[19] RD_M[19] VSS VSS VCC VCC RD[19] sky130_fd_sc_hd__inv_1
xRBUF[20] RD_M[20] VSS VSS VCC VCC RD[20] sky130_fd_sc_hd__inv_1
xRBUF[21] RD_M[21] VSS VSS VCC VCC RD[21] sky130_fd_sc_hd__inv_1
xRBUF[22] RD_M[22] VSS VSS VCC VCC RD[22] sky130_fd_sc_hd__inv_1
xRBUF[23] RD_M[23] VSS VSS VCC VCC RD[23] sky130_fd_sc_hd__inv_1
xRBUF[24] RD_M[24] VSS VSS VCC VCC RD[24] sky130_fd_sc_hd__inv_1
xRBUF[25] RD_M[25] VSS VSS VCC VCC RD[25] sky130_fd_sc_hd__inv_1
xRBUF[26] RD_M[26] VSS VSS VCC VCC RD[26] sky130_fd_sc_hd__inv_1
xRBUF[27] RD_M[27] VSS VSS VCC VCC RD[27] sky130_fd_sc_hd__inv_1
xRBUF[28] RD_M[28] VSS VSS VCC VCC RD[28] sky130_fd_sc_hd__inv_1
xRBUF[29] RD_M[29] VSS VSS VCC VCC RD[29] sky130_fd_sc_hd__inv_1
xRBUF[30] RD_M[30] VSS VSS VCC VCC RD[30] sky130_fd_sc_hd__inv_1
xRBUF[31] RD_M[31] VSS VSS VCC VCC RD[31] sky130_fd_sc_hd__inv_1
