* NGSPICE file created from rv_fetch.ext - technology: sky130A

.subckt rv_fetch
+ i_clk i_reset_n i_stall
+ i_pc_select i_ebreak
+ i_pc_target[1] i_pc_target[2] i_pc_target[3] i_pc_target[4] i_pc_target[5] i_pc_target[6] i_pc_target[7] i_pc_target[8] i_pc_target[9] i_pc_target[10] i_pc_target[11] i_pc_target[12] i_pc_target[13] i_pc_target[14] i_pc_target[15] 
+ i_pc_trap[1] i_pc_trap[2] i_pc_trap[3] i_pc_trap[4] i_pc_trap[5] i_pc_trap[6] i_pc_trap[7] i_pc_trap[8] i_pc_trap[9] i_pc_trap[10] i_pc_trap[11] i_pc_trap[12] i_pc_trap[13] i_pc_trap[14] i_pc_trap[15] 
+ i_ack o_cyc
+ i_instruction[0] i_instruction[1] i_instruction[2] i_instruction[3] i_instruction[4] i_instruction[5] i_instruction[6] i_instruction[7] i_instruction[8] i_instruction[9] i_instruction[10] i_instruction[11] i_instruction[12] i_instruction[13] i_instruction[14] i_instruction[15] i_instruction[16] i_instruction[17] i_instruction[18] i_instruction[19] i_instruction[20] i_instruction[21] i_instruction[22] i_instruction[23] i_instruction[24] i_instruction[25] i_instruction[26] i_instruction[27] i_instruction[28] i_instruction[29] i_instruction[30] i_instruction[31] 
+ o_addr[1] o_addr[2] o_addr[3] o_addr[4] o_addr[5] o_addr[6] o_addr[7] o_addr[8] o_addr[9] o_addr[10] o_addr[11] o_addr[12] o_addr[13] o_addr[14] o_addr[15] 
+ o_pc_change o_ready
+ o_pc[1] o_pc[2] o_pc[3] o_pc[4] o_pc[5] o_pc[6] o_pc[7] o_pc[8] o_pc[9] o_pc[10] o_pc[11] o_pc[12] o_pc[13] o_pc[14] o_pc[15] 
+ o_pc_next[1] o_pc_next[2] o_pc_next[3] o_pc_next[4] o_pc_next[5] o_pc_next[6] o_pc_next[7] o_pc_next[8] o_pc_next[9] o_pc_next[10] o_pc_next[11] o_pc_next[12] o_pc_next[13] o_pc_next[14] o_pc_next[15] 
+ o_instruction[0] o_instruction[1] o_instruction[2] o_instruction[3] o_instruction[4] o_instruction[5] o_instruction[6] o_instruction[7] o_instruction[8] o_instruction[9] o_instruction[10] o_instruction[11] o_instruction[12] o_instruction[13] o_instruction[14] o_instruction[15] o_instruction[16] o_instruction[17] o_instruction[18] o_instruction[19] o_instruction[20] o_instruction[21] o_instruction[22] o_instruction[23] o_instruction[24] o_instruction[25] o_instruction[26] o_instruction[27] o_instruction[28] o_instruction[29] o_instruction[30] o_instruction[31] 
+ vccd1 vssd1
X_0985_ _0059_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__clkbuf_1
X_0419_ _0072_ vssd1 vssd1 vccd1 vccd1 o_instruction[19] sky130_fd_sc_hd__buf_2
X_0770_ o_pc[5] _0287_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__and2_1
X_0968_ u_buf.data\[0\]\[21\] u_buf.latch_hi\[5\] _0045_ vssd1 vssd1 vccd1 vccd1 _0051_
+ sky130_fd_sc_hd__mux2_1
X_0899_ u_buf.is_head\[4\] _0378_ _0379_ u_buf.is_head\[2\] vssd1 vssd1 vccd1 vccd1
+ _0381_ sky130_fd_sc_hd__a22o_1
X_0822_ _0264_ _0339_ _0340_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__and3_1
X_0684_ i_instruction[15] _0223_ _0224_ u_buf.data\[0\]\[15\] vssd1 vssd1 vccd1 vccd1
+ _0230_ sky130_fd_sc_hd__a22o_1
X_0753_ o_pc[2] _0267_ o_pc[3] vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__a21o_1
X_1167_ clknet_4_10_0_i_clk o_pc_next[11] vssd1 vssd1 vccd1 vccd1 o_pc[11] sky130_fd_sc_hd__dfxtp_4
X_1098_ clknet_4_0_0_i_clk u_buf.g_data\[0\].d_next\[5\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_1021_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[27\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_0805_ o_pc[5] _0287_ _0324_ o_pc[9] vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__a31o_1
X_0736_ _0106_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__inv_2
X_0667_ i_instruction[8] _0209_ _0211_ u_buf.data\[0\]\[8\] vssd1 vssd1 vccd1 vccd1
+ _0220_ sky130_fd_sc_hd__a22o_1
X_0598_ u_buf.data\[1\]\[11\] _0178_ _0175_ i_instruction[11] _0179_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[11\] sky130_fd_sc_hd__a221o_1
X_0521_ u_buf.data\[3\]\[13\] _0129_ _0123_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__and3_1
X_0452_ u_buf.data\[0\]\[3\] u_buf.latch_hi\[3\] _0088_ vssd1 vssd1 vccd1 vccd1 _0090_
+ sky130_fd_sc_hd__mux2_1
X_1004_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[10\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_0719_ i_instruction[31] _0206_ _0210_ u_buf.data\[0\]\[31\] vssd1 vssd1 vccd1 vccd1
+ _0249_ sky130_fd_sc_hd__a22o_1
X_0435_ u_buf.data\[0\]\[27\] u_buf.data\[0\]\[11\] _0077_ vssd1 vssd1 vccd1 vccd1
+ _0081_ sky130_fd_sc_hd__mux2_1
X_0504_ u_buf.data\[2\]\[6\] _0109_ _0112_ i_instruction[6] _0122_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[6\] sky130_fd_sc_hd__a221o_1
X_0984_ u_buf.data\[0\]\[29\] u_buf.latch_hi\[13\] _0250_ vssd1 vssd1 vccd1 vccd1
+ _0059_ sky130_fd_sc_hd__mux2_1
X_0418_ u_buf.data\[0\]\[19\] u_buf.data\[0\]\[3\] _0068_ vssd1 vssd1 vccd1 vccd1
+ _0072_ sky130_fd_sc_hd__mux2_1
X_0967_ _0050_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__clkbuf_1
X_0898_ _0378_ _0379_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__nor2_1
X_0752_ o_pc[2] o_pc[3] _0267_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__nand3_1
X_0821_ o_pc[10] o_pc[11] _0325_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__nand3_1
X_0683_ u_buf.data\[1\]\[14\] _0222_ _0229_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[14\]
+ sky130_fd_sc_hd__a21o_1
X_1166_ clknet_4_10_0_i_clk o_pc_next[10] vssd1 vssd1 vccd1 vccd1 o_pc[10] sky130_fd_sc_hd__dfxtp_4
X_1097_ clknet_4_0_0_i_clk u_buf.g_data\[0\].d_next\[4\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_1020_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[26\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_0735_ _0263_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__buf_2
X_0804_ o_pc[5] o_pc[9] _0287_ _0324_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__and4_1
X_0666_ u_buf.data\[1\]\[7\] _0208_ _0219_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[7\]
+ sky130_fd_sc_hd__a21o_1
X_0597_ u_buf.data\[2\]\[11\] _0173_ _0176_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__and3_1
X_1149_ clknet_4_2_0_i_clk _0025_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[9\] sky130_fd_sc_hd__dfxtp_1
X_0520_ u_buf.data\[2\]\[12\] _0127_ _0128_ i_instruction[12] _0132_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[12\] sky130_fd_sc_hd__a221o_1
X_0451_ _0089_ vssd1 vssd1 vccd1 vccd1 o_instruction[2] sky130_fd_sc_hd__buf_2
X_1003_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[9\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_0718_ u_buf.data\[1\]\[30\] _0207_ _0248_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[30\]
+ sky130_fd_sc_hd__a21o_1
X_0649_ _0107_ _0205_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__nor2_2
Xclkbuf_4_15_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0434_ _0080_ vssd1 vssd1 vccd1 vccd1 o_instruction[26] sky130_fd_sc_hd__buf_2
X_0503_ u_buf.data\[3\]\[6\] _0113_ _0115_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__and3_1
X_0983_ _0058_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__clkbuf_1
X_0417_ _0071_ vssd1 vssd1 vccd1 vccd1 o_instruction[18] sky130_fd_sc_hd__buf_2
X_0966_ u_buf.data\[0\]\[20\] u_buf.latch_hi\[4\] _0045_ vssd1 vssd1 vccd1 vccd1 _0050_
+ sky130_fd_sc_hd__mux2_1
X_0897_ u_buf.i_push _0204_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__and2_1
X_0751_ _0255_ i_pc_trap[3] _0277_ _0065_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__o211a_1
X_0820_ o_pc[10] _0325_ o_pc[11] vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__a21o_1
X_0682_ i_instruction[14] _0223_ _0224_ u_buf.data\[0\]\[14\] vssd1 vssd1 vccd1 vccd1
+ _0229_ sky130_fd_sc_hd__a22o_1
X_1165_ clknet_4_10_0_i_clk o_pc_next[9] vssd1 vssd1 vccd1 vccd1 o_pc[9] sky130_fd_sc_hd__dfxtp_4
X_1096_ clknet_4_0_0_i_clk u_buf.g_data\[0\].d_next\[3\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_0949_ _0039_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__clkbuf_1
X_0734_ u_buf.first_half _0251_ _0262_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__and3b_1
X_0803_ o_pc[6] o_pc[7] o_pc[8] vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__and3_1
X_0665_ i_instruction[7] _0209_ _0211_ u_buf.data\[0\]\[7\] vssd1 vssd1 vccd1 vccd1
+ _0219_ sky130_fd_sc_hd__a22o_1
X_0596_ _0158_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__buf_2
X_1148_ clknet_4_0_0_i_clk _0024_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[8\] sky130_fd_sc_hd__dfxtp_1
X_1079_ clknet_4_12_0_i_clk u_buf.g_data\[1\].d_next\[19\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_0450_ u_buf.data\[0\]\[2\] u_buf.latch_hi\[2\] _0088_ vssd1 vssd1 vccd1 vccd1 _0089_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_11_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_1002_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[8\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_0648_ _0206_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__buf_2
X_0717_ i_instruction[30] _0206_ _0210_ u_buf.data\[0\]\[30\] vssd1 vssd1 vccd1 vccd1
+ _0248_ sky130_fd_sc_hd__a22o_1
X_0579_ u_buf.data\[2\]\[4\] _0161_ _0162_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__and3_1
X_0502_ u_buf.data\[2\]\[5\] _0109_ _0112_ i_instruction[5] _0121_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[5\] sky130_fd_sc_hd__a221o_1
X_0433_ u_buf.data\[0\]\[26\] u_buf.data\[0\]\[10\] _0077_ vssd1 vssd1 vccd1 vccd1
+ _0080_ sky130_fd_sc_hd__mux2_1
X_0982_ u_buf.data\[0\]\[28\] u_buf.latch_hi\[12\] _0250_ vssd1 vssd1 vccd1 vccd1
+ _0058_ sky130_fd_sc_hd__mux2_1
X_0416_ u_buf.data\[0\]\[18\] u_buf.data\[0\]\[2\] _0068_ vssd1 vssd1 vccd1 vccd1
+ _0071_ sky130_fd_sc_hd__mux2_1
X_0965_ _0049_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__clkbuf_1
X_0896_ u_buf.i_push _0204_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__nor2_1
X_0750_ _0270_ i_pc_target[3] _0275_ _0276_ i_ebreak vssd1 vssd1 vccd1 vccd1 _0277_
+ sky130_fd_sc_hd__a221o_1
X_0681_ u_buf.data\[1\]\[13\] _0222_ _0228_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[13\]
+ sky130_fd_sc_hd__a21o_1
X_1164_ clknet_4_10_0_i_clk o_pc_next[8] vssd1 vssd1 vccd1 vccd1 o_pc[8] sky130_fd_sc_hd__dfxtp_4
X_1095_ clknet_4_0_0_i_clk u_buf.g_data\[0\].d_next\[2\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_0948_ o_addr[13] _0354_ _0395_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__mux2_1
X_0879_ u_buf.data\[3\]\[18\] _0373_ _0374_ i_instruction[18] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[18\] sky130_fd_sc_hd__a22o_1
X_0802_ _0254_ i_pc_trap[9] _0321_ _0322_ i_reset_n vssd1 vssd1 vccd1 vccd1 _0323_
+ sky130_fd_sc_hd__o221a_1
X_0733_ _0250_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__inv_2
X_0664_ u_buf.data\[1\]\[6\] _0208_ _0218_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[6\]
+ sky130_fd_sc_hd__a21o_1
X_0595_ u_buf.data\[1\]\[10\] _0164_ _0175_ i_instruction[10] _0177_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[10\] sky130_fd_sc_hd__a221o_1
X_1078_ clknet_4_5_0_i_clk u_buf.g_data\[1\].d_next\[18\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_1147_ clknet_4_0_0_i_clk _0023_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[7\] sky130_fd_sc_hd__dfxtp_1
X_1001_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[7\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_0578_ u_buf.data\[1\]\[3\] _0164_ _0160_ i_instruction[3] _0167_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[3\] sky130_fd_sc_hd__a221o_1
X_0647_ _0207_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__buf_2
X_0716_ u_buf.data\[1\]\[29\] _0235_ _0247_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[29\]
+ sky130_fd_sc_hd__a21o_1
X_0432_ _0079_ vssd1 vssd1 vccd1 vccd1 o_instruction[25] sky130_fd_sc_hd__buf_2
X_0501_ u_buf.data\[3\]\[5\] _0113_ _0115_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_9_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0981_ _0057_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__clkbuf_1
X_0415_ _0070_ vssd1 vssd1 vccd1 vccd1 o_instruction[17] sky130_fd_sc_hd__buf_2
X_0964_ u_buf.data\[0\]\[19\] u_buf.latch_hi\[3\] _0045_ vssd1 vssd1 vccd1 vccd1 _0049_
+ sky130_fd_sc_hd__mux2_1
X_0895_ i_reset_n _0063_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__nand2_2
X_0680_ i_instruction[13] _0223_ _0224_ u_buf.data\[0\]\[13\] vssd1 vssd1 vccd1 vccd1
+ _0228_ sky130_fd_sc_hd__a22o_1
X_1163_ clknet_4_10_0_i_clk o_pc_next[7] vssd1 vssd1 vccd1 vccd1 o_pc[7] sky130_fd_sc_hd__dfxtp_4
X_1094_ clknet_4_3_0_i_clk u_buf.g_data\[0\].d_next\[1\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_0947_ o_addr[12] _0391_ _0037_ _0038_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a22o_1
X_0878_ u_buf.data\[3\]\[17\] _0373_ _0374_ i_instruction[17] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[17\] sky130_fd_sc_hd__a22o_1
X_0801_ _0270_ i_pc_target[9] _0258_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__a21o_1
X_0732_ u_buf.data\[0\]\[0\] u_buf.data\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__nand2_1
X_0663_ i_instruction[6] _0209_ _0211_ u_buf.data\[0\]\[6\] vssd1 vssd1 vccd1 vccd1
+ _0218_ sky130_fd_sc_hd__a22o_1
X_0594_ u_buf.data\[2\]\[10\] _0173_ _0176_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__and3_1
X_1146_ clknet_4_0_0_i_clk _0022_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[6\] sky130_fd_sc_hd__dfxtp_1
X_1077_ clknet_4_13_0_i_clk u_buf.g_data\[1\].d_next\[17\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_1000_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[6\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_0715_ i_instruction[29] _0236_ _0237_ u_buf.data\[0\]\[29\] vssd1 vssd1 vccd1 vccd1
+ _0247_ sky130_fd_sc_hd__a22o_1
X_0646_ _0204_ _0206_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__nor2_1
X_0577_ u_buf.data\[2\]\[3\] _0161_ _0162_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_5_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_1129_ clknet_4_11_0_i_clk _0005_ vssd1 vssd1 vccd1 vccd1 o_addr[5] sky130_fd_sc_hd__dfxtp_2
X_0431_ u_buf.data\[0\]\[25\] u_buf.data\[0\]\[9\] _0077_ vssd1 vssd1 vccd1 vccd1
+ _0079_ sky130_fd_sc_hd__mux2_1
X_0500_ u_buf.data\[2\]\[4\] _0109_ _0112_ i_instruction[4] _0120_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[4\] sky130_fd_sc_hd__a221o_1
X_0629_ u_buf.data\[2\]\[25\] _0187_ _0190_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__and3_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_0980_ u_buf.data\[0\]\[27\] u_buf.latch_hi\[11\] _0250_ vssd1 vssd1 vccd1 vccd1
+ _0057_ sky130_fd_sc_hd__mux2_1
X_0414_ u_buf.data\[0\]\[17\] u_buf.data\[0\]\[1\] _0068_ vssd1 vssd1 vccd1 vccd1
+ _0070_ sky130_fd_sc_hd__mux2_1
X_0963_ _0048_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__clkbuf_1
X_0894_ u_buf.data\[3\]\[31\] _0369_ _0371_ i_instruction[31] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[31\] sky130_fd_sc_hd__a22o_1
X_1162_ clknet_4_10_0_i_clk o_pc_next[6] vssd1 vssd1 vccd1 vccd1 o_pc[6] sky130_fd_sc_hd__dfxtp_4
X_1093_ clknet_4_2_0_i_clk u_buf.g_data\[0\].d_next\[0\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_0877_ u_buf.data\[3\]\[16\] _0373_ _0374_ i_instruction[16] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[16\] sky130_fd_sc_hd__a22o_1
X_0946_ _0346_ _0391_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__nor2_1
X_0731_ _0255_ i_pc_trap[1] _0259_ _0065_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__o211a_1
X_0800_ _0270_ _0319_ _0320_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__nor3b_1
X_0662_ u_buf.data\[1\]\[5\] _0208_ _0217_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[5\]
+ sky130_fd_sc_hd__a21o_1
X_0593_ _0157_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_2
X_1145_ clknet_4_0_0_i_clk _0021_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[5\] sky130_fd_sc_hd__dfxtp_1
X_1076_ clknet_4_5_0_i_clk u_buf.g_data\[1\].d_next\[16\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_1_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0929_ o_addr[6] _0301_ _0395_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__mux2_1
X_0645_ u_buf.is_head\[1\] _0107_ _0205_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__a21o_1
X_0714_ u_buf.data\[1\]\[28\] _0235_ _0246_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[28\]
+ sky130_fd_sc_hd__a21o_1
X_0576_ u_buf.data\[1\]\[2\] _0164_ _0160_ i_instruction[2] _0166_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[2\] sky130_fd_sc_hd__a221o_1
X_1128_ clknet_4_8_0_i_clk _0004_ vssd1 vssd1 vccd1 vccd1 o_addr[4] sky130_fd_sc_hd__dfxtp_4
X_1059_ clknet_4_11_0_i_clk u_buf.g_data\[1\].h_next vssd1 vssd1 vccd1 vccd1 u_buf.is_head\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_0430_ _0078_ vssd1 vssd1 vccd1 vccd1 o_instruction[24] sky130_fd_sc_hd__buf_2
X_0628_ u_buf.data\[1\]\[24\] _0192_ _0189_ i_instruction[24] _0196_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[24\] sky130_fd_sc_hd__a221o_1
X_0559_ u_buf.data\[3\]\[30\] _0110_ _0114_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__and3_1
X_0413_ _0069_ vssd1 vssd1 vccd1 vccd1 o_instruction[16] sky130_fd_sc_hd__buf_2
X_0962_ u_buf.data\[0\]\[18\] u_buf.latch_hi\[2\] _0045_ vssd1 vssd1 vccd1 vccd1 _0048_
+ sky130_fd_sc_hd__mux2_1
X_0893_ u_buf.data\[3\]\[30\] _0369_ _0371_ i_instruction[30] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[30\] sky130_fd_sc_hd__a22o_1
X_1161_ clknet_4_10_0_i_clk o_pc_next[5] vssd1 vssd1 vccd1 vccd1 o_pc[5] sky130_fd_sc_hd__dfxtp_4
X_1092_ clknet_4_9_0_i_clk u_buf.g_data\[0\].h_next vssd1 vssd1 vccd1 vccd1 u_buf.is_head\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_0876_ u_buf.data\[3\]\[15\] _0373_ _0374_ i_instruction[15] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[15\] sky130_fd_sc_hd__a22o_1
X_0945_ _0257_ _0036_ _0347_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__o21ai_1
X_0730_ _0257_ i_pc_target[1] _0258_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__a21o_1
X_0661_ i_instruction[5] _0209_ _0211_ u_buf.data\[0\]\[5\] vssd1 vssd1 vccd1 vccd1
+ _0217_ sky130_fd_sc_hd__a22o_1
X_0592_ _0159_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__buf_2
X_1075_ clknet_4_7_0_i_clk u_buf.g_data\[1\].d_next\[15\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_1144_ clknet_4_0_0_i_clk _0020_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[4\] sky130_fd_sc_hd__dfxtp_1
X_0928_ _0397_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__clkbuf_1
X_0859_ u_buf.data\[3\]\[0\] _0370_ _0372_ i_instruction[0] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[0\] sky130_fd_sc_hd__a22o_1
X_0644_ u_buf.i_push u_buf.is_head\[0\] vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__and2_1
X_0713_ i_instruction[28] _0236_ _0237_ u_buf.data\[0\]\[28\] vssd1 vssd1 vccd1 vccd1
+ _0246_ sky130_fd_sc_hd__a22o_1
X_0575_ u_buf.data\[2\]\[2\] _0161_ _0162_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__and3_1
X_1127_ clknet_4_8_0_i_clk _0003_ vssd1 vssd1 vccd1 vccd1 o_addr[3] sky130_fd_sc_hd__dfxtp_4
X_1058_ clknet_4_6_0_i_clk u_buf.g_data\[2\].d_next\[31\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_0558_ u_buf.data\[2\]\[29\] _0141_ _0142_ i_instruction[29] _0153_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[29\] sky130_fd_sc_hd__a221o_1
X_0627_ u_buf.data\[2\]\[24\] _0187_ _0190_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__and3_1
X_0489_ _0107_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__buf_2
X_0412_ u_buf.data\[0\]\[16\] u_buf.data\[0\]\[0\] _0068_ vssd1 vssd1 vccd1 vccd1
+ _0069_ sky130_fd_sc_hd__mux2_1
X_0961_ _0047_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__clkbuf_1
X_0892_ u_buf.data\[3\]\[29\] _0375_ _0376_ i_instruction[29] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[29\] sky130_fd_sc_hd__a22o_1
X_1160_ clknet_4_10_0_i_clk o_pc_next[4] vssd1 vssd1 vccd1 vccd1 o_pc[4] sky130_fd_sc_hd__dfxtp_4
X_1091_ clknet_4_9_0_i_clk u_buf.g_data\[1\].d_next\[31\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_0944_ o_addr[12] _0335_ _0349_ _0319_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__a2bb2o_1
X_0875_ u_buf.data\[3\]\[14\] _0373_ _0374_ i_instruction[14] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[14\] sky130_fd_sc_hd__a22o_1
X_0660_ u_buf.data\[1\]\[4\] _0208_ _0216_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[4\]
+ sky130_fd_sc_hd__a21o_1
X_0591_ u_buf.data\[1\]\[9\] _0164_ _0160_ i_instruction[9] _0174_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[9\] sky130_fd_sc_hd__a221o_1
X_1143_ clknet_4_0_0_i_clk _0019_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[3\] sky130_fd_sc_hd__dfxtp_1
X_1074_ clknet_4_7_0_i_clk u_buf.g_data\[1\].d_next\[14\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_0927_ o_addr[5] _0294_ _0395_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__mux2_1
X_0789_ _0310_ _0311_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__nor2_1
X_0858_ _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__buf_2
X_0643_ u_buf.hi_valid _0106_ _0103_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__a21o_1
X_0574_ u_buf.data\[1\]\[1\] _0164_ _0160_ i_instruction[1] _0165_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[1\] sky130_fd_sc_hd__a221o_1
X_0712_ u_buf.data\[1\]\[27\] _0235_ _0245_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[27\]
+ sky130_fd_sc_hd__a21o_1
X_1126_ clknet_4_8_0_i_clk _0002_ vssd1 vssd1 vccd1 vccd1 o_addr[2] sky130_fd_sc_hd__dfxtp_4
X_1057_ clknet_4_12_0_i_clk u_buf.g_data\[2\].d_next\[30\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_0557_ u_buf.data\[3\]\[29\] _0143_ _0114_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__and3_1
X_0626_ u_buf.data\[1\]\[23\] _0192_ _0189_ i_instruction[23] _0195_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[23\] sky130_fd_sc_hd__a221o_1
X_0488_ _0110_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__clkbuf_2
X_1109_ clknet_4_5_0_i_clk u_buf.g_data\[0\].d_next\[16\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_0411_ _0067_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkbuf_4
X_0609_ u_buf.data\[2\]\[17\] _0173_ _0176_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__and3_1
X_0960_ u_buf.data\[0\]\[17\] u_buf.latch_hi\[1\] _0045_ vssd1 vssd1 vccd1 vccd1 _0047_
+ sky130_fd_sc_hd__mux2_1
X_0891_ u_buf.data\[3\]\[28\] _0375_ _0376_ i_instruction[28] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[28\] sky130_fd_sc_hd__a22o_1
X_1090_ clknet_4_12_0_i_clk u_buf.g_data\[1\].d_next\[30\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_0874_ u_buf.data\[3\]\[13\] _0373_ _0374_ i_instruction[13] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[13\] sky130_fd_sc_hd__a22o_1
X_0943_ _0035_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__clkbuf_1
X_0590_ u_buf.data\[2\]\[9\] _0173_ _0162_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__and3_1
X_1142_ clknet_4_0_0_i_clk _0018_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[2\] sky130_fd_sc_hd__dfxtp_1
X_1073_ clknet_4_7_0_i_clk u_buf.g_data\[1\].d_next\[13\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_0926_ _0396_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__clkbuf_1
X_0857_ u_buf.is_head\[4\] _0114_ _0368_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__a21o_1
X_0788_ o_pc[7] _0302_ _0264_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__o21ai_1
X_0711_ i_instruction[27] _0236_ _0237_ u_buf.data\[0\]\[27\] vssd1 vssd1 vccd1 vccd1
+ _0245_ sky130_fd_sc_hd__a22o_1
X_0573_ u_buf.data\[2\]\[1\] _0161_ _0162_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__and3_1
X_0642_ u_buf.data\[1\]\[31\] _0158_ _0159_ i_instruction[31] _0203_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[31\] sky130_fd_sc_hd__a221o_1
X_1125_ clknet_4_14_0_i_clk _0001_ vssd1 vssd1 vccd1 vccd1 o_addr[1] sky130_fd_sc_hd__dfxtp_2
X_1056_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[29\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_0909_ u_buf.hi_valid u_buf.is_head\[0\] _0068_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__and3b_1
X_0625_ u_buf.data\[2\]\[23\] _0187_ _0190_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__and3_1
X_0556_ u_buf.data\[2\]\[28\] _0141_ _0142_ i_instruction[28] _0152_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[28\] sky130_fd_sc_hd__a221o_1
X_0487_ _0111_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__buf_2
X_1039_ clknet_4_5_0_i_clk u_buf.g_data\[2\].d_next\[12\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_1108_ clknet_4_6_0_i_clk u_buf.g_data\[0\].d_next\[15\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_0410_ o_pc[1] vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__buf_2
X_0608_ u_buf.data\[1\]\[16\] _0178_ _0175_ i_instruction[16] _0184_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[16\] sky130_fd_sc_hd__a221o_1
X_0539_ u_buf.data\[3\]\[20\] _0143_ _0137_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__and3_1
X_0890_ u_buf.data\[3\]\[27\] _0375_ _0376_ i_instruction[27] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[27\] sky130_fd_sc_hd__a22o_1
X_0873_ u_buf.data\[3\]\[12\] _0373_ _0374_ i_instruction[12] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[12\] sky130_fd_sc_hd__a22o_1
X_0942_ o_addr[11] _0338_ _0395_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__mux2_1
X_1141_ clknet_4_2_0_i_clk _0017_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[1\] sky130_fd_sc_hd__dfxtp_1
X_1072_ clknet_4_5_0_i_clk u_buf.g_data\[1\].d_next\[12\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_0787_ o_pc[7] _0302_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__and2_1
X_0925_ o_addr[4] _0286_ _0395_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__mux2_1
X_0856_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__buf_2
X_0641_ u_buf.data\[2\]\[31\] _0115_ _0157_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__and3_1
X_0710_ u_buf.data\[1\]\[26\] _0235_ _0244_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[26\]
+ sky130_fd_sc_hd__a21o_1
X_0572_ _0158_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__buf_2
X_1055_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[28\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_1124_ clknet_4_9_0_i_clk u_buf.g_data\[0\].d_next\[31\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_0839_ o_pc[13] _0343_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__nand2_1
X_0908_ u_buf.is_head\[0\] u_buf.first_half vssd1 vssd1 vccd1 vccd1 o_ready sky130_fd_sc_hd__nor2_4
X_0624_ u_buf.data\[1\]\[22\] _0192_ _0189_ i_instruction[22] _0194_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[22\] sky130_fd_sc_hd__a221o_1
X_0555_ u_buf.data\[3\]\[28\] _0143_ _0114_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__and3_1
X_0486_ _0110_ _0108_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__nor2_1
X_1107_ clknet_4_6_0_i_clk u_buf.g_data\[0\].d_next\[14\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_1038_ clknet_4_5_0_i_clk u_buf.g_data\[2\].d_next\[11\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_0538_ _0110_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__clkbuf_2
X_0607_ u_buf.data\[2\]\[16\] _0173_ _0176_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__and3_1
X_0469_ _0098_ vssd1 vssd1 vccd1 vccd1 o_instruction[11] sky130_fd_sc_hd__buf_2
X_0941_ _0034_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__clkbuf_1
X_0872_ u_buf.data\[3\]\[11\] _0373_ _0374_ i_instruction[11] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[11\] sky130_fd_sc_hd__a22o_1
X_1140_ clknet_4_0_0_i_clk _0016_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[0\] sky130_fd_sc_hd__dfxtp_1
X_1071_ clknet_4_5_0_i_clk u_buf.g_data\[1\].d_next\[11\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_0924_ _0391_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__inv_2
X_0786_ _0255_ i_pc_trap[7] _0308_ _0065_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__o211a_1
X_0855_ _0114_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__nor2_2
X_0571_ i_instruction[0] _0160_ _0163_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[1\].d_next\[0\]
+ sky130_fd_sc_hd__a21o_1
X_0640_ u_buf.data\[1\]\[30\] _0192_ _0159_ i_instruction[30] _0202_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[30\] sky130_fd_sc_hd__a221o_1
X_1123_ clknet_4_12_0_i_clk u_buf.g_data\[0\].d_next\[30\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_1054_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[27\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_0907_ _0386_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].h_next sky130_fd_sc_hd__clkbuf_1
X_0838_ o_pc[13] _0343_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__or2_1
X_0769_ _0254_ i_pc_trap[5] _0292_ _0293_ i_reset_n vssd1 vssd1 vccd1 vccd1 _0294_
+ sky130_fd_sc_hd__o221a_1
X_0623_ u_buf.data\[2\]\[22\] _0187_ _0190_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__and3_1
X_0554_ u_buf.data\[2\]\[27\] _0141_ _0142_ i_instruction[27] _0151_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[27\] sky130_fd_sc_hd__a221o_1
X_0485_ u_buf.is_head\[3\] _0105_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__nor2_2
X_1106_ clknet_4_7_0_i_clk u_buf.g_data\[0\].d_next\[13\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_1037_ clknet_4_5_0_i_clk u_buf.g_data\[2\].d_next\[10\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_14_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0537_ _0111_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__buf_2
X_0606_ u_buf.data\[1\]\[15\] _0178_ _0175_ i_instruction[15] _0183_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[15\] sky130_fd_sc_hd__a221o_1
X_0468_ u_buf.data\[0\]\[11\] u_buf.latch_hi\[11\] _0088_ vssd1 vssd1 vccd1 vccd1
+ _0098_ sky130_fd_sc_hd__mux2_1
X_0940_ o_addr[10] _0331_ _0395_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__mux2_1
X_0871_ u_buf.data\[3\]\[10\] _0373_ _0374_ i_instruction[10] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[10\] sky130_fd_sc_hd__a22o_1
X_1070_ clknet_4_4_0_i_clk u_buf.g_data\[1\].d_next\[10\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_0923_ _0394_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__clkbuf_1
X_0854_ u_buf.is_head\[3\] u_buf.i_push _0104_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__and3_1
X_0785_ _0256_ i_pc_target[7] _0305_ _0307_ i_ebreak vssd1 vssd1 vccd1 vccd1 _0308_
+ sky130_fd_sc_hd__a221o_1
X_0570_ u_buf.data\[2\]\[0\] _0161_ _0162_ _0158_ u_buf.data\[1\]\[0\] vssd1 vssd1
+ vccd1 vccd1 _0163_ sky130_fd_sc_hd__a32o_1
X_1122_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[29\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_1053_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[26\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_0906_ _0251_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__and2_1
X_0837_ _0254_ i_pc_trap[13] _0352_ _0353_ i_reset_n vssd1 vssd1 vccd1 vccd1 _0354_
+ sky130_fd_sc_hd__o221a_1
X_0768_ _0270_ i_pc_target[5] _0258_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__a21o_1
X_0699_ i_instruction[21] _0236_ _0237_ u_buf.data\[0\]\[21\] vssd1 vssd1 vccd1 vccd1
+ _0239_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_10_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0553_ u_buf.data\[3\]\[27\] _0143_ _0114_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__and3_1
X_0484_ _0108_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__buf_2
X_0622_ u_buf.data\[1\]\[21\] _0192_ _0189_ i_instruction[21] _0193_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[21\] sky130_fd_sc_hd__a221o_1
X_1105_ clknet_4_4_0_i_clk u_buf.g_data\[0\].d_next\[12\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_1036_ clknet_4_6_0_i_clk u_buf.g_data\[2\].d_next\[9\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_0605_ u_buf.data\[2\]\[15\] _0173_ _0176_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__and3_1
X_0536_ _0108_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__buf_2
X_0467_ _0097_ vssd1 vssd1 vccd1 vccd1 o_instruction[10] sky130_fd_sc_hd__buf_2
X_1019_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[25\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_0519_ u_buf.data\[3\]\[12\] _0129_ _0123_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__and3_1
X_0870_ _0371_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__buf_2
X_0999_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[5\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_0853_ o_pc[15] _0252_ _0365_ _0264_ _0367_ vssd1 vssd1 vccd1 vccd1 o_pc_next[15]
+ sky130_fd_sc_hd__a221o_4
X_0922_ _0278_ o_addr[3] _0391_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__mux2_1
X_0784_ _0256_ _0306_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__nor2_1
X_1052_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[25\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_1121_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[28\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_0767_ _0257_ _0290_ _0291_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__nor3_1
X_0905_ u_buf.is_head\[2\] _0378_ _0380_ u_buf.is_head\[1\] _0205_ vssd1 vssd1 vccd1
+ vccd1 _0385_ sky130_fd_sc_hd__a221o_1
X_0836_ _0270_ i_pc_target[13] _0258_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__a21o_1
X_0698_ u_buf.data\[1\]\[20\] _0235_ _0238_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[20\]
+ sky130_fd_sc_hd__a21o_1
X_0621_ u_buf.data\[2\]\[21\] _0187_ _0190_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__and3_1
X_0552_ u_buf.data\[2\]\[26\] _0141_ _0142_ i_instruction[26] _0150_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[26\] sky130_fd_sc_hd__a221o_1
X_0483_ _0105_ _0107_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__nor2_2
X_1035_ clknet_4_3_0_i_clk u_buf.g_data\[2\].d_next\[8\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_1104_ clknet_4_4_0_i_clk u_buf.g_data\[0\].d_next\[11\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_0819_ _0254_ i_pc_trap[11] _0336_ _0337_ i_reset_n vssd1 vssd1 vccd1 vccd1 _0338_
+ sky130_fd_sc_hd__o221a_1
X_0604_ u_buf.data\[1\]\[14\] _0178_ _0175_ i_instruction[14] _0182_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[14\] sky130_fd_sc_hd__a221o_1
X_0535_ u_buf.data\[2\]\[19\] _0127_ _0128_ i_instruction[19] _0140_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[19\] sky130_fd_sc_hd__a221o_1
X_0466_ u_buf.data\[0\]\[10\] u_buf.latch_hi\[10\] _0088_ vssd1 vssd1 vccd1 vccd1
+ _0097_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_8_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_1018_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[24\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_0518_ u_buf.data\[2\]\[11\] _0127_ _0128_ i_instruction[11] _0131_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[11\] sky130_fd_sc_hd__a221o_1
X_0449_ _0067_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__clkbuf_4
X_0998_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[4\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_0921_ _0393_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__clkbuf_1
X_0852_ _0255_ i_pc_trap[15] _0366_ _0065_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__o211a_1
X_0783_ o_addr[6] o_addr[7] _0290_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__and3_1
X_1051_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[24\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_1120_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[27\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_0904_ _0377_ _0384_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[1\].h_next sky130_fd_sc_hd__nor2_1
X_0766_ o_addr[5] _0283_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__nor2_1
X_0835_ _0257_ _0350_ _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__nor3_1
X_0697_ i_instruction[20] _0236_ _0237_ u_buf.data\[0\]\[20\] vssd1 vssd1 vccd1 vccd1
+ _0238_ sky130_fd_sc_hd__a22o_1
X_0551_ u_buf.data\[3\]\[26\] _0143_ _0137_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__and3_1
X_0620_ _0158_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__buf_2
X_0482_ u_buf.hi_valid _0106_ _0103_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__a21oi_4
X_1034_ clknet_4_1_0_i_clk u_buf.g_data\[2\].d_next\[7\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_1103_ clknet_4_5_0_i_clk u_buf.g_data\[0\].d_next\[10\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_4_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0749_ o_addr[2] o_addr[3] _0256_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__o21ba_1
X_0818_ _0270_ i_pc_target[11] _0258_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__a21o_1
X_0534_ u_buf.data\[3\]\[19\] _0129_ _0137_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__and3_1
X_0603_ u_buf.data\[2\]\[14\] _0173_ _0176_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__and3_1
X_0465_ _0096_ vssd1 vssd1 vccd1 vccd1 o_instruction[9] sky130_fd_sc_hd__buf_2
X_1017_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[23\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_0517_ u_buf.data\[3\]\[11\] _0129_ _0123_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__and3_1
X_0448_ _0087_ vssd1 vssd1 vccd1 vccd1 o_instruction[1] sky130_fd_sc_hd__buf_2
X_0997_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[3\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_0920_ _0273_ _0392_ _0391_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__mux2_1
X_0782_ o_addr[6] _0290_ o_addr[7] vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__a21o_1
X_0851_ _0257_ i_pc_target[15] _0258_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__a21o_1
X_1050_ clknet_4_15_0_i_clk u_buf.g_data\[2\].d_next\[23\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_0834_ o_addr[13] _0319_ _0349_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__and3_1
X_0903_ u_buf.is_head\[2\] _0380_ _0383_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__a21oi_1
X_0765_ o_addr[2] o_addr[3] o_addr[4] o_addr[5] vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__and4_2
X_0696_ _0210_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__buf_2
Xclkbuf_4_0_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0550_ u_buf.data\[2\]\[25\] _0141_ _0142_ i_instruction[25] _0149_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[25\] sky130_fd_sc_hd__a221o_1
X_0481_ u_buf.latch_hi\[0\] u_buf.latch_hi\[1\] _0067_ vssd1 vssd1 vccd1 vccd1 _0106_
+ sky130_fd_sc_hd__a21boi_4
X_1102_ clknet_4_3_0_i_clk u_buf.g_data\[0\].d_next\[9\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_1033_ clknet_4_1_0_i_clk u_buf.g_data\[2\].d_next\[6\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_0817_ _0257_ _0334_ _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__nor3_1
X_0748_ o_addr[2] o_addr[3] vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__nand2_1
X_0679_ u_buf.data\[1\]\[12\] _0222_ _0227_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[12\]
+ sky130_fd_sc_hd__a21o_1
X_0533_ u_buf.data\[2\]\[18\] _0127_ _0128_ i_instruction[18] _0139_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[18\] sky130_fd_sc_hd__a221o_1
X_0602_ u_buf.data\[1\]\[13\] _0178_ _0175_ i_instruction[13] _0181_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[13\] sky130_fd_sc_hd__a221o_1
X_0464_ u_buf.data\[0\]\[9\] u_buf.latch_hi\[9\] _0088_ vssd1 vssd1 vccd1 vccd1 _0096_
+ sky130_fd_sc_hd__mux2_1
X_1016_ clknet_4_13_0_i_clk u_buf.g_data\[3\].d_next\[22\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_0516_ u_buf.data\[2\]\[10\] _0127_ _0128_ i_instruction[10] _0130_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[10\] sky130_fd_sc_hd__a221o_1
X_0447_ u_buf.data\[0\]\[1\] u_buf.latch_hi\[1\] _0077_ vssd1 vssd1 vccd1 vccd1 _0087_
+ sky130_fd_sc_hd__mux2_1
X_0996_ clknet_4_4_0_i_clk u_buf.g_data\[3\].d_next\[2\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_0850_ o_pc[15] _0362_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__xor2_1
X_0781_ o_pc[6] _0253_ _0301_ o_pc_change _0304_ vssd1 vssd1 vccd1 vccd1 o_pc_next[6]
+ sky130_fd_sc_hd__a221o_4
X_0979_ _0056_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__clkbuf_1
X_0902_ u_buf.is_head\[3\] _0378_ _0379_ u_buf.is_head\[1\] vssd1 vssd1 vccd1 vccd1
+ _0383_ sky130_fd_sc_hd__a22o_1
X_0833_ _0319_ _0349_ o_addr[13] vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__a21oi_1
X_0764_ o_pc[4] _0253_ _0286_ o_pc_change _0289_ vssd1 vssd1 vccd1 vccd1 o_pc_next[4]
+ sky130_fd_sc_hd__a221o_4
X_0695_ _0206_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__buf_2
X_0480_ u_buf.i_push u_buf.is_head\[2\] _0104_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__and3_1
X_1101_ clknet_4_2_0_i_clk u_buf.g_data\[0\].d_next\[8\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_1032_ clknet_4_1_0_i_clk u_buf.g_data\[2\].d_next\[5\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_0747_ o_pc[2] _0251_ _0268_ _0274_ vssd1 vssd1 vccd1 vccd1 o_pc_next[2] sky130_fd_sc_hd__a31o_4
X_0816_ o_addr[10] o_addr[11] _0319_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__and3_1
X_0678_ i_instruction[12] _0223_ _0224_ u_buf.data\[0\]\[12\] vssd1 vssd1 vccd1 vccd1
+ _0227_ sky130_fd_sc_hd__a22o_1
X_0601_ u_buf.data\[2\]\[13\] _0173_ _0176_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__and3_1
X_0532_ u_buf.data\[3\]\[18\] _0129_ _0137_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__and3_1
X_0463_ _0095_ vssd1 vssd1 vccd1 vccd1 o_instruction[8] sky130_fd_sc_hd__buf_2
X_1015_ clknet_4_13_0_i_clk u_buf.g_data\[3\].d_next\[21\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_0515_ u_buf.data\[3\]\[10\] _0129_ _0123_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__and3_1
X_0446_ _0086_ vssd1 vssd1 vccd1 vccd1 o_instruction[0] sky130_fd_sc_hd__buf_2
X_0995_ clknet_4_6_0_i_clk u_buf.g_data\[3\].d_next\[1\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_0429_ u_buf.data\[0\]\[24\] u_buf.data\[0\]\[8\] _0077_ vssd1 vssd1 vccd1 vccd1
+ _0078_ sky130_fd_sc_hd__mux2_1
X_0780_ _0302_ _0303_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__nor2_1
X_0978_ u_buf.data\[0\]\[26\] u_buf.latch_hi\[10\] _0250_ vssd1 vssd1 vccd1 vccd1
+ _0056_ sky130_fd_sc_hd__mux2_1
X_0763_ _0287_ _0288_ _0263_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__and3b_1
X_0832_ o_addr[10] o_addr[11] o_addr[12] vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__and3_1
X_0901_ _0377_ _0382_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[2\].h_next sky130_fd_sc_hd__nor2_1
X_0694_ _0207_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__buf_2
X_1100_ clknet_4_2_0_i_clk u_buf.g_data\[0\].d_next\[7\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_1031_ clknet_4_4_0_i_clk u_buf.g_data\[2\].d_next\[4\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_0746_ _0269_ _0264_ _0267_ _0273_ _0064_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__a32o_1
X_0815_ o_addr[10] _0319_ o_addr[11] vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__a21oi_1
X_0677_ u_buf.data\[1\]\[11\] _0222_ _0226_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[11\]
+ sky130_fd_sc_hd__a21o_1
X_0531_ u_buf.data\[2\]\[17\] _0127_ _0128_ i_instruction[17] _0138_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[17\] sky130_fd_sc_hd__a221o_1
X_0600_ u_buf.data\[1\]\[12\] _0178_ _0175_ i_instruction[12] _0180_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[12\] sky130_fd_sc_hd__a221o_1
X_0462_ u_buf.data\[0\]\[8\] u_buf.latch_hi\[8\] _0088_ vssd1 vssd1 vccd1 vccd1 _0095_
+ sky130_fd_sc_hd__mux2_1
X_1014_ clknet_4_13_0_i_clk u_buf.g_data\[3\].d_next\[20\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_0729_ i_ebreak vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__buf_2
X_0514_ _0110_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__clkbuf_2
X_0445_ u_buf.data\[0\]\[0\] u_buf.latch_hi\[0\] _0077_ vssd1 vssd1 vccd1 vccd1 _0086_
+ sky130_fd_sc_hd__mux2_1
X_0994_ clknet_4_6_0_i_clk u_buf.g_data\[3\].d_next\[0\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_0428_ _0067_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__clkbuf_4
X_0977_ _0055_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__clkbuf_1
X_0900_ u_buf.is_head\[3\] _0380_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__a21oi_1
X_0831_ o_pc[12] _0253_ _0345_ _0348_ vssd1 vssd1 vccd1 vccd1 o_pc_next[12] sky130_fd_sc_hd__a211o_4
X_0762_ o_pc[2] o_pc[3] _0267_ o_pc[4] vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__a31o_1
X_0693_ u_buf.data\[1\]\[19\] _0222_ _0234_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[19\]
+ sky130_fd_sc_hd__a21o_1
X_1030_ clknet_4_1_0_i_clk u_buf.g_data\[2\].d_next\[3\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_0814_ o_pc[10] _0253_ _0331_ o_pc_change _0333_ vssd1 vssd1 vccd1 vccd1 o_pc_next[10]
+ sky130_fd_sc_hd__a221o_4
X_0745_ _0254_ i_pc_trap[2] _0272_ i_reset_n vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__o211a_1
X_0676_ i_instruction[11] _0223_ _0224_ u_buf.data\[0\]\[11\] vssd1 vssd1 vccd1 vccd1
+ _0226_ sky130_fd_sc_hd__a22o_1
X_1159_ clknet_4_8_0_i_clk o_pc_next[3] vssd1 vssd1 vccd1 vccd1 o_pc[3] sky130_fd_sc_hd__dfxtp_4
X_0530_ u_buf.data\[3\]\[17\] _0129_ _0137_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__and3_1
X_0461_ _0094_ vssd1 vssd1 vccd1 vccd1 o_instruction[7] sky130_fd_sc_hd__buf_2
X_1013_ clknet_4_13_0_i_clk u_buf.g_data\[3\].d_next\[19\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_0728_ _0256_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__buf_2
X_0659_ i_instruction[4] _0209_ _0211_ u_buf.data\[0\]\[4\] vssd1 vssd1 vccd1 vccd1
+ _0216_ sky130_fd_sc_hd__a22o_1
X_0513_ _0111_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__buf_2
X_0444_ _0085_ vssd1 vssd1 vccd1 vccd1 o_instruction[31] sky130_fd_sc_hd__buf_2
X_0993_ clknet_4_9_0_i_clk u_buf.g_data\[3\].h_next vssd1 vssd1 vccd1 vccd1 u_buf.is_head\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_0427_ _0076_ vssd1 vssd1 vccd1 vccd1 o_instruction[23] sky130_fd_sc_hd__buf_2
X_0976_ u_buf.data\[0\]\[25\] u_buf.latch_hi\[9\] _0045_ vssd1 vssd1 vccd1 vccd1 _0055_
+ sky130_fd_sc_hd__mux2_1
X_0830_ _0346_ _0347_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__nor2_1
X_0761_ o_pc[2] o_pc[3] o_pc[4] _0267_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__and4_1
X_0692_ i_instruction[19] _0223_ _0224_ u_buf.data\[0\]\[19\] vssd1 vssd1 vccd1 vccd1
+ _0234_ sky130_fd_sc_hd__a22o_1
X_0959_ _0046_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__clkbuf_1
X_0813_ o_pc[10] _0325_ _0332_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__o21a_1
X_0744_ _0270_ i_pc_target[2] _0271_ _0258_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__a211o_1
X_0675_ u_buf.data\[1\]\[10\] _0222_ _0225_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[10\]
+ sky130_fd_sc_hd__a21o_1
X_1158_ clknet_4_8_0_i_clk o_pc_next[2] vssd1 vssd1 vccd1 vccd1 o_pc[2] sky130_fd_sc_hd__dfxtp_4
X_1089_ clknet_4_14_0_i_clk u_buf.g_data\[1\].d_next\[29\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_0460_ u_buf.data\[0\]\[7\] u_buf.latch_hi\[7\] _0088_ vssd1 vssd1 vccd1 vccd1 _0094_
+ sky130_fd_sc_hd__mux2_1
X_1012_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[18\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_0727_ i_pc_select vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__buf_2
X_0658_ u_buf.data\[1\]\[3\] _0208_ _0215_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[3\]
+ sky130_fd_sc_hd__a21o_1
X_0589_ _0114_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_2
X_0512_ _0108_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__buf_2
X_0443_ u_buf.data\[0\]\[31\] u_buf.data\[0\]\[15\] _0077_ vssd1 vssd1 vccd1 vccd1
+ _0085_ sky130_fd_sc_hd__mux2_1
X_0992_ clknet_4_9_0_i_clk u_buf.is_head_next_0 vssd1 vssd1 vccd1 vccd1 u_buf.is_head\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_0426_ u_buf.data\[0\]\[23\] u_buf.data\[0\]\[7\] _0068_ vssd1 vssd1 vccd1 vccd1
+ _0076_ sky130_fd_sc_hd__mux2_1
X_0975_ _0054_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__clkbuf_1
X_0409_ _0066_ vssd1 vssd1 vccd1 vccd1 push_next sky130_fd_sc_hd__clkbuf_1
X_0760_ _0255_ i_pc_trap[4] _0285_ _0065_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__o211a_1
X_0691_ u_buf.data\[1\]\[18\] _0222_ _0233_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[18\]
+ sky130_fd_sc_hd__a21o_1
X_0889_ u_buf.data\[3\]\[26\] _0375_ _0376_ i_instruction[26] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[26\] sky130_fd_sc_hd__a22o_1
X_0958_ u_buf.data\[0\]\[16\] u_buf.latch_hi\[0\] _0045_ vssd1 vssd1 vccd1 vccd1 _0046_
+ sky130_fd_sc_hd__mux2_1
X_0812_ o_pc[10] _0325_ _0263_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__a21boi_1
X_0743_ _0256_ o_addr[2] vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__nor2_1
X_0674_ i_instruction[10] _0223_ _0224_ u_buf.data\[0\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _0225_ sky130_fd_sc_hd__a22o_1
X_1157_ clknet_4_8_0_i_clk o_pc_next[1] vssd1 vssd1 vccd1 vccd1 o_pc[1] sky130_fd_sc_hd__dfxtp_2
X_1088_ clknet_4_14_0_i_clk u_buf.g_data\[1\].d_next\[28\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_1011_ clknet_4_7_0_i_clk u_buf.g_data\[3\].d_next\[17\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_0726_ _0254_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__buf_2
X_0657_ i_instruction[3] _0209_ _0211_ u_buf.data\[0\]\[3\] vssd1 vssd1 vccd1 vccd1
+ _0215_ sky130_fd_sc_hd__a22o_1
X_0588_ u_buf.data\[1\]\[8\] _0164_ _0160_ i_instruction[8] _0172_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[8\] sky130_fd_sc_hd__a221o_1
X_0511_ u_buf.data\[2\]\[9\] _0109_ _0112_ i_instruction[9] _0126_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[9\] sky130_fd_sc_hd__a221o_1
Xclkbuf_4_13_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0442_ _0084_ vssd1 vssd1 vccd1 vccd1 o_instruction[30] sky130_fd_sc_hd__buf_2
X_0709_ i_instruction[26] _0236_ _0237_ u_buf.data\[0\]\[26\] vssd1 vssd1 vccd1 vccd1
+ _0244_ sky130_fd_sc_hd__a22o_1
X_0991_ _0377_ _0062_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__nor2_1
X_0425_ _0075_ vssd1 vssd1 vccd1 vccd1 o_instruction[22] sky130_fd_sc_hd__buf_2
X_0974_ u_buf.data\[0\]\[24\] u_buf.latch_hi\[8\] _0045_ vssd1 vssd1 vccd1 vccd1 _0054_
+ sky130_fd_sc_hd__mux2_1
X_0408_ _0065_ i_ack _0063_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__and3_1
X_0690_ i_instruction[18] _0223_ _0224_ u_buf.data\[0\]\[18\] vssd1 vssd1 vccd1 vccd1
+ _0233_ sky130_fd_sc_hd__a22o_1
X_1173_ clknet_4_9_0_i_clk push_next vssd1 vssd1 vccd1 vccd1 u_buf.i_push sky130_fd_sc_hd__dfxtp_2
X_0888_ u_buf.data\[3\]\[25\] _0375_ _0376_ i_instruction[25] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[25\] sky130_fd_sc_hd__a22o_1
X_0957_ _0250_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__clkbuf_4
X_0811_ _0254_ i_pc_trap[10] _0330_ i_reset_n vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__o211a_1
X_0742_ _0256_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__buf_2
X_0673_ _0210_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__buf_2
X_1156_ clknet_4_8_0_i_clk _0000_ vssd1 vssd1 vccd1 vccd1 u_buf.first_half sky130_fd_sc_hd__dfxtp_1
X_1087_ clknet_4_14_0_i_clk u_buf.g_data\[1\].d_next\[27\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_1010_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[16\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_0725_ i_ebreak vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkinv_2
X_0656_ u_buf.data\[1\]\[2\] _0208_ _0214_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[2\]
+ sky130_fd_sc_hd__a21o_1
X_0587_ u_buf.data\[2\]\[8\] _0161_ _0162_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__and3_1
X_1139_ clknet_4_11_0_i_clk _0015_ vssd1 vssd1 vccd1 vccd1 o_addr[15] sky130_fd_sc_hd__dfxtp_4
X_0510_ u_buf.data\[3\]\[9\] _0113_ _0123_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__and3_1
X_0441_ u_buf.data\[0\]\[30\] u_buf.data\[0\]\[14\] _0077_ vssd1 vssd1 vccd1 vccd1
+ _0084_ sky130_fd_sc_hd__mux2_1
X_0639_ u_buf.data\[2\]\[30\] _0115_ _0157_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__and3_1
X_0708_ u_buf.data\[1\]\[25\] _0235_ _0243_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[25\]
+ sky130_fd_sc_hd__a21o_1
X_0990_ u_buf.i_push _0262_ u_buf.hi_valid vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__a21oi_1
X_0424_ u_buf.data\[0\]\[22\] u_buf.data\[0\]\[6\] _0068_ vssd1 vssd1 vccd1 vccd1
+ _0075_ sky130_fd_sc_hd__mux2_1
X_0973_ _0053_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__clkbuf_1
X_0407_ i_reset_n vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__buf_2
X_1172_ clknet_4_8_0_i_clk _0032_ vssd1 vssd1 vccd1 vccd1 u_buf.hi_valid sky130_fd_sc_hd__dfxtp_1
X_0956_ o_addr[15] _0391_ _0043_ _0044_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a22o_1
X_0887_ u_buf.data\[3\]\[24\] _0375_ _0376_ i_instruction[24] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[24\] sky130_fd_sc_hd__a22o_1
X_0810_ _0256_ i_pc_target[10] _0328_ _0329_ i_ebreak vssd1 vssd1 vccd1 vccd1 _0330_
+ sky130_fd_sc_hd__a221o_1
X_0741_ o_pc[2] vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__inv_2
X_0672_ _0206_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__buf_2
X_1155_ clknet_4_8_0_i_clk _0031_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[15\] sky130_fd_sc_hd__dfxtp_1
X_1086_ clknet_4_15_0_i_clk u_buf.g_data\[1\].d_next\[26\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_0939_ _0033_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__clkbuf_1
X_0724_ _0252_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__buf_4
X_0655_ i_instruction[2] _0209_ _0211_ u_buf.data\[0\]\[2\] vssd1 vssd1 vccd1 vccd1
+ _0214_ sky130_fd_sc_hd__a22o_1
X_0586_ u_buf.data\[1\]\[7\] _0164_ _0160_ i_instruction[7] _0171_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[7\] sky130_fd_sc_hd__a221o_1
X_1069_ clknet_4_3_0_i_clk u_buf.g_data\[1\].d_next\[9\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_1138_ clknet_4_11_0_i_clk _0014_ vssd1 vssd1 vccd1 vccd1 o_addr[14] sky130_fd_sc_hd__dfxtp_4
X_0440_ _0083_ vssd1 vssd1 vccd1 vccd1 o_instruction[29] sky130_fd_sc_hd__buf_2
X_0707_ i_instruction[25] _0236_ _0237_ u_buf.data\[0\]\[25\] vssd1 vssd1 vccd1 vccd1
+ _0243_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_7_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0569_ _0157_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_2
X_0638_ u_buf.data\[1\]\[29\] _0192_ _0189_ i_instruction[29] _0201_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[29\] sky130_fd_sc_hd__a221o_1
X_0423_ _0074_ vssd1 vssd1 vccd1 vccd1 o_instruction[21] sky130_fd_sc_hd__buf_2
X_0972_ u_buf.data\[0\]\[23\] u_buf.latch_hi\[7\] _0045_ vssd1 vssd1 vccd1 vccd1 _0053_
+ sky130_fd_sc_hd__mux2_1
X_0406_ _0064_ vssd1 vssd1 vccd1 vccd1 o_pc_change sky130_fd_sc_hd__buf_6
X_1171_ clknet_4_10_0_i_clk o_pc_next[15] vssd1 vssd1 vccd1 vccd1 o_pc[15] sky130_fd_sc_hd__dfxtp_4
X_0886_ u_buf.data\[3\]\[23\] _0375_ _0376_ i_instruction[23] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[23\] sky130_fd_sc_hd__a22o_1
X_0955_ _0255_ i_pc_trap[15] _0395_ _0065_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__o211a_1
X_0740_ u_buf.first_half _0250_ _0267_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__or3b_1
X_0671_ _0207_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__buf_2
X_1154_ clknet_4_2_0_i_clk _0030_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[14\] sky130_fd_sc_hd__dfxtp_1
X_1085_ clknet_4_14_0_i_clk u_buf.g_data\[1\].d_next\[25\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_0869_ _0369_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__buf_2
X_0938_ o_addr[9] _0323_ _0395_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__mux2_1
X_0723_ u_buf.first_half _0250_ _0251_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__o21a_2
X_0654_ u_buf.data\[1\]\[1\] _0208_ _0213_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[1\]
+ sky130_fd_sc_hd__a21o_1
X_0585_ u_buf.data\[2\]\[7\] _0161_ _0162_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_3_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_1137_ clknet_4_11_0_i_clk _0013_ vssd1 vssd1 vccd1 vccd1 o_addr[13] sky130_fd_sc_hd__dfxtp_4
X_1068_ clknet_4_3_0_i_clk u_buf.g_data\[1\].d_next\[8\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_0706_ u_buf.data\[1\]\[24\] _0235_ _0242_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[24\]
+ sky130_fd_sc_hd__a21o_1
X_0568_ _0107_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_2
X_0499_ u_buf.data\[3\]\[4\] _0113_ _0115_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__and3_1
X_0637_ u_buf.data\[2\]\[29\] _0115_ _0190_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__and3_1
X_0422_ u_buf.data\[0\]\[21\] u_buf.data\[0\]\[5\] _0068_ vssd1 vssd1 vccd1 vccd1
+ _0074_ sky130_fd_sc_hd__mux2_1
X_0971_ _0052_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__clkbuf_1
X_0405_ _0063_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__inv_2
X_1170_ clknet_4_10_0_i_clk o_pc_next[14] vssd1 vssd1 vccd1 vccd1 o_pc[14] sky130_fd_sc_hd__dfxtp_4
X_0885_ u_buf.data\[3\]\[22\] _0375_ _0376_ i_instruction[22] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[22\] sky130_fd_sc_hd__a22o_1
X_0954_ _0041_ _0042_ _0366_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__a21o_1
X_0670_ u_buf.data\[1\]\[9\] _0208_ _0221_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[9\]
+ sky130_fd_sc_hd__a21o_1
X_1153_ clknet_4_2_0_i_clk _0029_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[13\] sky130_fd_sc_hd__dfxtp_1
X_1084_ clknet_4_14_0_i_clk u_buf.g_data\[1\].d_next\[24\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_0799_ o_addr[6] _0290_ _0317_ o_addr[9] vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__a31o_1
X_0937_ o_addr[8] _0391_ _0402_ _0403_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__a22o_1
X_0868_ u_buf.data\[3\]\[9\] _0370_ _0372_ i_instruction[9] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[9\] sky130_fd_sc_hd__a22o_1
X_0722_ i_reset_n _0063_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__and2_1
X_0653_ i_instruction[1] _0209_ _0211_ u_buf.data\[0\]\[1\] vssd1 vssd1 vccd1 vccd1
+ _0213_ sky130_fd_sc_hd__a22o_1
X_0584_ u_buf.data\[1\]\[6\] _0164_ _0160_ i_instruction[6] _0170_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[6\] sky130_fd_sc_hd__a221o_1
X_1136_ clknet_4_11_0_i_clk _0012_ vssd1 vssd1 vccd1 vccd1 o_addr[12] sky130_fd_sc_hd__dfxtp_2
X_1067_ clknet_4_1_0_i_clk u_buf.g_data\[1\].d_next\[7\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_0705_ i_instruction[24] _0236_ _0237_ u_buf.data\[0\]\[24\] vssd1 vssd1 vccd1 vccd1
+ _0242_ sky130_fd_sc_hd__a22o_1
X_0636_ u_buf.data\[1\]\[28\] _0192_ _0189_ i_instruction[28] _0200_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[28\] sky130_fd_sc_hd__a221o_1
X_0567_ _0159_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__buf_2
X_0498_ u_buf.data\[2\]\[3\] _0109_ _0112_ i_instruction[3] _0119_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[3\] sky130_fd_sc_hd__a221o_1
X_1119_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[26\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_0421_ _0073_ vssd1 vssd1 vccd1 vccd1 o_instruction[20] sky130_fd_sc_hd__buf_2
X_0619_ u_buf.data\[1\]\[20\] _0178_ _0189_ i_instruction[20] _0191_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[20\] sky130_fd_sc_hd__a221o_1
X_0970_ u_buf.data\[0\]\[22\] u_buf.latch_hi\[6\] _0045_ vssd1 vssd1 vccd1 vccd1 _0052_
+ sky130_fd_sc_hd__mux2_1
X_0404_ i_ebreak i_pc_select vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__nor2_1
X_0884_ u_buf.data\[3\]\[21\] _0375_ _0376_ i_instruction[21] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[21\] sky130_fd_sc_hd__a22o_1
X_0953_ o_addr[14] o_addr[15] _0351_ _0257_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__a31oi_1
X_1152_ clknet_4_2_0_i_clk _0028_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[12\] sky130_fd_sc_hd__dfxtp_1
X_1083_ clknet_4_15_0_i_clk u_buf.g_data\[1\].d_next\[23\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_0936_ _0314_ _0391_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__nor2_1
X_0798_ _0318_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__clkbuf_2
X_0867_ u_buf.data\[3\]\[8\] _0370_ _0372_ i_instruction[8] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[8\] sky130_fd_sc_hd__a22o_1
X_0721_ _0103_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__clkbuf_4
X_0652_ u_buf.data\[1\]\[0\] _0208_ _0212_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[0\]
+ sky130_fd_sc_hd__a21o_1
X_0583_ u_buf.data\[2\]\[6\] _0161_ _0162_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__and3_1
X_1135_ clknet_4_10_0_i_clk _0011_ vssd1 vssd1 vccd1 vccd1 o_addr[11] sky130_fd_sc_hd__dfxtp_4
X_1066_ clknet_4_3_0_i_clk u_buf.g_data\[1\].d_next\[6\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_0919_ _0255_ i_pc_trap[2] _0272_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__o21ai_1
X_0566_ _0157_ _0158_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__nor2_1
X_0704_ u_buf.data\[1\]\[23\] _0235_ _0241_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[23\]
+ sky130_fd_sc_hd__a21o_1
X_0635_ u_buf.data\[2\]\[28\] _0187_ _0190_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__and3_1
X_0497_ u_buf.data\[3\]\[3\] _0113_ _0115_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__and3_1
X_1049_ clknet_4_13_0_i_clk u_buf.g_data\[2\].d_next\[22\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_1118_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[25\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_0420_ u_buf.data\[0\]\[20\] u_buf.data\[0\]\[4\] _0068_ vssd1 vssd1 vccd1 vccd1
+ _0073_ sky130_fd_sc_hd__mux2_1
X_0549_ u_buf.data\[3\]\[25\] _0143_ _0137_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__and3_1
X_0618_ u_buf.data\[2\]\[20\] _0187_ _0190_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__and3_1
X_0952_ o_addr[14] _0351_ o_addr[15] vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__a21o_1
X_0883_ u_buf.data\[3\]\[20\] _0375_ _0376_ i_instruction[20] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[20\] sky130_fd_sc_hd__a22o_1
X_1151_ clknet_4_2_0_i_clk _0027_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[11\] sky130_fd_sc_hd__dfxtp_1
X_1082_ clknet_4_13_0_i_clk u_buf.g_data\[1\].d_next\[22\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_0935_ _0257_ _0401_ _0315_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__o21ai_1
X_0866_ u_buf.data\[3\]\[7\] _0370_ _0372_ i_instruction[7] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[7\] sky130_fd_sc_hd__a22o_1
X_0797_ o_addr[6] o_addr[9] _0290_ _0317_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__and4_1
X_0720_ u_buf.data\[1\]\[31\] _0207_ _0249_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[31\]
+ sky130_fd_sc_hd__a21o_1
X_0582_ u_buf.data\[1\]\[5\] _0164_ _0160_ i_instruction[5] _0169_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[5\] sky130_fd_sc_hd__a221o_1
X_0651_ i_instruction[0] _0209_ _0211_ u_buf.data\[0\]\[0\] vssd1 vssd1 vccd1 vccd1
+ _0212_ sky130_fd_sc_hd__a22o_1
X_1134_ clknet_4_11_0_i_clk _0010_ vssd1 vssd1 vccd1 vccd1 o_addr[10] sky130_fd_sc_hd__dfxtp_4
X_1065_ clknet_4_1_0_i_clk u_buf.g_data\[1\].d_next\[5\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_0849_ o_pc[14] _0252_ _0361_ _0064_ _0364_ vssd1 vssd1 vccd1 vccd1 o_pc_next[14]
+ sky130_fd_sc_hd__a221o_4
X_0918_ o_addr[1] _0391_ _0260_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a21o_1
X_0703_ i_instruction[23] _0236_ _0237_ u_buf.data\[0\]\[23\] vssd1 vssd1 vccd1 vccd1
+ _0241_ sky130_fd_sc_hd__a22o_1
X_0565_ _0107_ _0156_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__nor2_2
X_0496_ u_buf.data\[2\]\[2\] _0109_ _0112_ i_instruction[2] _0118_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[2\] sky130_fd_sc_hd__a221o_1
X_0634_ u_buf.data\[1\]\[27\] _0192_ _0189_ i_instruction[27] _0199_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[27\] sky130_fd_sc_hd__a221o_1
X_1117_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[24\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_1048_ clknet_4_13_0_i_clk u_buf.g_data\[2\].d_next\[21\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_0548_ u_buf.data\[2\]\[24\] _0141_ _0142_ i_instruction[24] _0148_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[24\] sky130_fd_sc_hd__a221o_1
X_0479_ _0067_ _0103_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__or2_1
X_0617_ _0157_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_2
X_0882_ _0371_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__buf_2
X_0951_ _0040_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__clkbuf_1
X_1150_ clknet_4_2_0_i_clk _0026_ vssd1 vssd1 vccd1 vccd1 u_buf.latch_hi\[10\] sky130_fd_sc_hd__dfxtp_1
X_1081_ clknet_4_13_0_i_clk u_buf.g_data\[1\].d_next\[21\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_0934_ o_addr[6] _0290_ _0317_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__a31o_1
X_0865_ u_buf.data\[3\]\[6\] _0370_ _0372_ i_instruction[6] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[6\] sky130_fd_sc_hd__a22o_1
X_0796_ o_addr[7] o_addr[8] vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__and2_1
X_0650_ _0210_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__buf_2
X_0581_ u_buf.data\[2\]\[5\] _0161_ _0162_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__and3_1
X_1064_ clknet_4_1_0_i_clk u_buf.g_data\[1\].d_next\[4\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_1133_ clknet_4_11_0_i_clk _0009_ vssd1 vssd1 vccd1 vccd1 o_addr[9] sky130_fd_sc_hd__dfxtp_2
X_0848_ _0362_ _0263_ _0363_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__and3b_1
X_0779_ o_pc[6] _0295_ _0264_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__o21ai_1
X_0917_ i_ack o_cyc _0377_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__a21oi_4
X_0702_ u_buf.data\[1\]\[22\] _0235_ _0240_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[22\]
+ sky130_fd_sc_hd__a21o_1
X_0633_ u_buf.data\[2\]\[27\] _0187_ _0190_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__and3_1
X_0564_ u_buf.is_head\[2\] _0156_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__nor2_2
X_0495_ u_buf.data\[3\]\[2\] _0113_ _0115_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__and3_1
X_1047_ clknet_4_13_0_i_clk u_buf.g_data\[2\].d_next\[20\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_1116_ clknet_4_14_0_i_clk u_buf.g_data\[0\].d_next\[23\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_0616_ _0159_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__buf_2
X_0547_ u_buf.data\[3\]\[24\] _0143_ _0137_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__and3_1
X_0478_ u_buf.is_head\[0\] i_stall vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__or2_2
X_0881_ _0369_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__buf_2
X_0950_ o_addr[14] _0361_ _0395_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__mux2_1
X_1080_ clknet_4_13_0_i_clk u_buf.g_data\[1\].d_next\[20\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_0795_ o_pc[8] _0253_ _0313_ _0264_ _0316_ vssd1 vssd1 vccd1 vccd1 o_pc_next[8] sky130_fd_sc_hd__a221o_4
X_0933_ o_addr[8] _0306_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__nor2_1
X_0864_ u_buf.data\[3\]\[5\] _0370_ _0372_ i_instruction[5] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[5\] sky130_fd_sc_hd__a22o_1
X_0580_ u_buf.data\[1\]\[4\] _0164_ _0160_ i_instruction[4] _0168_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[4\] sky130_fd_sc_hd__a221o_1
X_1063_ clknet_4_1_0_i_clk u_buf.g_data\[1\].d_next\[3\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1132_ clknet_4_11_0_i_clk _0008_ vssd1 vssd1 vccd1 vccd1 o_addr[8] sky130_fd_sc_hd__dfxtp_4
X_0916_ _0390_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[3\].h_next sky130_fd_sc_hd__clkbuf_1
X_0847_ o_pc[13] _0343_ o_pc[14] vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__a21o_1
X_0778_ o_pc[5] o_pc[6] _0287_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__and3_1
X_0563_ u_buf.i_push u_buf.is_head\[1\] _0104_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__and3_1
X_0701_ i_instruction[22] _0236_ _0237_ u_buf.data\[0\]\[22\] vssd1 vssd1 vccd1 vccd1
+ _0240_ sky130_fd_sc_hd__a22o_1
X_0632_ u_buf.data\[1\]\[26\] _0192_ _0189_ i_instruction[26] _0198_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[26\] sky130_fd_sc_hd__a221o_1
X_0494_ u_buf.data\[2\]\[1\] _0109_ _0112_ i_instruction[1] _0117_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[1\] sky130_fd_sc_hd__a221o_1
X_1046_ clknet_4_13_0_i_clk u_buf.g_data\[2\].d_next\[19\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_1115_ clknet_4_12_0_i_clk u_buf.g_data\[0\].d_next\[22\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_0546_ u_buf.data\[2\]\[23\] _0141_ _0142_ i_instruction[23] _0147_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[23\] sky130_fd_sc_hd__a221o_1
X_0615_ u_buf.data\[1\]\[19\] _0178_ _0175_ i_instruction[19] _0188_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[19\] sky130_fd_sc_hd__a221o_1
X_0477_ _0102_ vssd1 vssd1 vccd1 vccd1 o_instruction[15] sky130_fd_sc_hd__buf_2
X_1029_ clknet_4_1_0_i_clk u_buf.g_data\[2\].d_next\[2\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_0529_ _0107_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__clkbuf_2
X_0880_ u_buf.data\[3\]\[19\] _0373_ _0374_ i_instruction[19] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[19\] sky130_fd_sc_hd__a22o_1
X_0932_ _0399_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__clkbuf_1
X_0794_ _0314_ _0315_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__nor2_1
X_0863_ u_buf.data\[3\]\[4\] _0370_ _0372_ i_instruction[4] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[4\] sky130_fd_sc_hd__a22o_1
X_1131_ clknet_4_11_0_i_clk _0007_ vssd1 vssd1 vccd1 vccd1 o_addr[7] sky130_fd_sc_hd__dfxtp_4
X_1062_ clknet_4_1_0_i_clk u_buf.g_data\[1\].d_next\[2\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_0915_ _0251_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__and2_1
X_0846_ o_pc[13] o_pc[14] _0343_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__and3_1
X_0777_ _0255_ i_pc_trap[6] _0300_ _0065_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__o211a_1
X_0700_ u_buf.data\[1\]\[21\] _0235_ _0239_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[21\]
+ sky130_fd_sc_hd__a21o_1
X_0562_ u_buf.data\[2\]\[31\] _0108_ _0111_ i_instruction[31] _0155_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[31\] sky130_fd_sc_hd__a221o_1
X_0631_ u_buf.data\[2\]\[26\] _0187_ _0190_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__and3_1
X_0493_ u_buf.data\[3\]\[1\] _0113_ _0115_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__and3_1
X_1114_ clknet_4_12_0_i_clk u_buf.g_data\[0\].d_next\[21\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_1045_ clknet_4_7_0_i_clk u_buf.g_data\[2\].d_next\[18\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_0829_ _0257_ i_pc_target[12] _0258_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_4_12_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0545_ u_buf.data\[3\]\[23\] _0143_ _0137_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__and3_1
X_0476_ u_buf.data\[0\]\[15\] u_buf.latch_hi\[15\] _0067_ vssd1 vssd1 vccd1 vccd1
+ _0102_ sky130_fd_sc_hd__mux2_1
X_0614_ u_buf.data\[2\]\[19\] _0187_ _0176_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__and3_1
X_1028_ clknet_4_3_0_i_clk u_buf.g_data\[2\].d_next\[1\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_0528_ u_buf.data\[2\]\[16\] _0127_ _0128_ i_instruction[16] _0136_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[16\] sky130_fd_sc_hd__a221o_1
X_0459_ _0093_ vssd1 vssd1 vccd1 vccd1 o_instruction[6] sky130_fd_sc_hd__buf_2
X_0931_ o_addr[7] _0309_ _0395_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__mux2_1
X_0862_ u_buf.data\[3\]\[3\] _0370_ _0372_ i_instruction[3] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[3\] sky130_fd_sc_hd__a22o_1
X_0793_ _0257_ i_pc_target[8] _0258_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a21oi_1
X_1130_ clknet_4_10_0_i_clk _0006_ vssd1 vssd1 vccd1 vccd1 o_addr[6] sky130_fd_sc_hd__dfxtp_4
X_1061_ clknet_4_3_0_i_clk u_buf.g_data\[1\].d_next\[1\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_0914_ u_buf.is_head\[3\] _0379_ _0380_ u_buf.is_head\[4\] vssd1 vssd1 vccd1 vccd1
+ _0389_ sky130_fd_sc_hd__a22o_1
X_0845_ _0254_ i_pc_trap[14] _0359_ _0360_ i_reset_n vssd1 vssd1 vccd1 vccd1 _0361_
+ sky130_fd_sc_hd__o221a_1
X_0776_ _0270_ i_pc_target[6] _0298_ _0299_ i_ebreak vssd1 vssd1 vccd1 vccd1 _0300_
+ sky130_fd_sc_hd__a221o_1
X_0492_ u_buf.data\[2\]\[0\] _0109_ _0112_ i_instruction[0] _0116_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[0\] sky130_fd_sc_hd__a221o_1
X_0561_ u_buf.data\[3\]\[31\] _0110_ _0114_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__and3_1
X_0630_ u_buf.data\[1\]\[25\] _0192_ _0189_ i_instruction[25] _0197_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[25\] sky130_fd_sc_hd__a221o_1
X_1044_ clknet_4_7_0_i_clk u_buf.g_data\[2\].d_next\[17\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_1113_ clknet_4_12_0_i_clk u_buf.g_data\[0\].d_next\[20\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_0828_ _0255_ i_pc_trap[12] _0065_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__o21ai_1
X_0759_ _0270_ i_pc_target[4] _0282_ _0284_ i_ebreak vssd1 vssd1 vccd1 vccd1 _0285_
+ sky130_fd_sc_hd__a221o_1
X_0613_ _0114_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__clkbuf_2
X_0544_ u_buf.data\[2\]\[22\] _0141_ _0142_ i_instruction[22] _0146_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[22\] sky130_fd_sc_hd__a221o_1
X_0475_ _0101_ vssd1 vssd1 vccd1 vccd1 o_instruction[14] sky130_fd_sc_hd__buf_2
X_1027_ clknet_4_3_0_i_clk u_buf.g_data\[2\].d_next\[0\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_0527_ u_buf.data\[3\]\[16\] _0129_ _0123_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__and3_1
X_0458_ u_buf.data\[0\]\[6\] u_buf.latch_hi\[6\] _0088_ vssd1 vssd1 vccd1 vccd1 _0093_
+ sky130_fd_sc_hd__mux2_1
X_0930_ _0398_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__clkbuf_1
X_0792_ _0255_ i_pc_trap[8] _0065_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__o21ai_1
X_0861_ u_buf.data\[3\]\[2\] _0370_ _0372_ i_instruction[2] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[2\] sky130_fd_sc_hd__a22o_1
X_1060_ clknet_4_3_0_i_clk u_buf.g_data\[1\].d_next\[0\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_0913_ u_buf.is_head\[3\] u_buf.i_push _0103_ u_buf.is_head\[4\] vssd1 vssd1 vccd1
+ vccd1 o_cyc sky130_fd_sc_hd__a31oi_4
X_0775_ o_addr[6] _0290_ _0256_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__o21ba_1
X_0844_ _0270_ i_pc_target[14] _0258_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__a21o_1
X_0491_ u_buf.data\[3\]\[0\] _0113_ _0115_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__and3_1
X_0560_ u_buf.data\[2\]\[30\] _0108_ _0111_ i_instruction[30] _0154_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[30\] sky130_fd_sc_hd__a221o_1
X_1043_ clknet_4_5_0_i_clk u_buf.g_data\[2\].d_next\[16\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_1112_ clknet_4_6_0_i_clk u_buf.g_data\[0\].d_next\[19\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_0827_ _0343_ _0344_ _0264_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__and3b_1
X_0758_ _0256_ _0283_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__nor2_1
X_0689_ u_buf.data\[1\]\[17\] _0222_ _0232_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[17\]
+ sky130_fd_sc_hd__a21o_1
X_0612_ u_buf.data\[1\]\[18\] _0178_ _0175_ i_instruction[18] _0186_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[18\] sky130_fd_sc_hd__a221o_1
X_0543_ u_buf.data\[3\]\[22\] _0143_ _0137_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__and3_1
X_0474_ u_buf.data\[0\]\[14\] u_buf.latch_hi\[14\] _0067_ vssd1 vssd1 vccd1 vccd1
+ _0101_ sky130_fd_sc_hd__mux2_1
X_1026_ clknet_4_9_0_i_clk u_buf.g_data\[2\].h_next vssd1 vssd1 vccd1 vccd1 u_buf.is_head\[3\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_4_6_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0526_ u_buf.data\[2\]\[15\] _0127_ _0128_ i_instruction[15] _0135_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[15\] sky130_fd_sc_hd__a221o_1
X_0457_ _0092_ vssd1 vssd1 vccd1 vccd1 o_instruction[5] sky130_fd_sc_hd__buf_2
X_1009_ clknet_4_7_0_i_clk u_buf.g_data\[3\].d_next\[15\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_0509_ u_buf.data\[2\]\[8\] _0109_ _0112_ i_instruction[8] _0125_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[8\] sky130_fd_sc_hd__a221o_1
X_0791_ o_pc[8] _0310_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__xor2_1
X_0860_ u_buf.data\[3\]\[1\] _0370_ _0372_ i_instruction[1] vssd1 vssd1 vccd1 vccd1
+ u_buf.g_data\[3\].d_next\[1\] sky130_fd_sc_hd__a22o_1
X_0989_ _0061_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__clkbuf_1
X_0912_ u_buf.i_push _0388_ _0251_ vssd1 vssd1 vccd1 vccd1 u_buf.is_head_next_0 sky130_fd_sc_hd__o21ai_1
X_0774_ o_addr[6] _0290_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__nand2_1
X_0843_ o_addr[14] _0351_ _0358_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__o21ba_1
X_0490_ _0114_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__clkbuf_2
X_1042_ clknet_4_7_0_i_clk u_buf.g_data\[2\].d_next\[15\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_1111_ clknet_4_7_0_i_clk u_buf.g_data\[0\].d_next\[18\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_0826_ o_pc[10] o_pc[11] _0325_ o_pc[12] vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__a31o_1
X_0757_ o_addr[2] o_addr[3] o_addr[4] vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_2_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0688_ i_instruction[17] _0223_ _0224_ u_buf.data\[0\]\[17\] vssd1 vssd1 vccd1 vccd1
+ _0232_ sky130_fd_sc_hd__a22o_1
X_0611_ u_buf.data\[2\]\[18\] _0173_ _0176_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__and3_1
X_0542_ u_buf.data\[2\]\[21\] _0141_ _0142_ i_instruction[21] _0145_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[21\] sky130_fd_sc_hd__a221o_1
X_0473_ _0100_ vssd1 vssd1 vccd1 vccd1 o_instruction[13] sky130_fd_sc_hd__buf_2
X_1025_ clknet_4_6_0_i_clk u_buf.g_data\[3\].d_next\[31\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_0809_ o_addr[10] _0319_ i_pc_select vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__o21ba_1
X_0525_ u_buf.data\[3\]\[15\] _0129_ _0123_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__and3_1
X_0456_ u_buf.data\[0\]\[5\] u_buf.latch_hi\[5\] _0088_ vssd1 vssd1 vccd1 vccd1 _0092_
+ sky130_fd_sc_hd__mux2_1
X_1008_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[14\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_0439_ u_buf.data\[0\]\[29\] u_buf.data\[0\]\[13\] _0077_ vssd1 vssd1 vccd1 vccd1
+ _0083_ sky130_fd_sc_hd__mux2_1
X_0508_ u_buf.data\[3\]\[8\] _0113_ _0123_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__and3_1
X_0790_ o_pc[7] _0253_ _0309_ o_pc_change _0312_ vssd1 vssd1 vccd1 vccd1 o_pc_next[7]
+ sky130_fd_sc_hd__a221o_4
X_0988_ u_buf.data\[0\]\[31\] u_buf.latch_hi\[15\] _0250_ vssd1 vssd1 vccd1 vccd1
+ _0061_ sky130_fd_sc_hd__mux2_1
X_0911_ u_buf.is_head\[1\] _0161_ u_buf.is_head\[0\] vssd1 vssd1 vccd1 vccd1 _0388_
+ sky130_fd_sc_hd__a21oi_1
X_0842_ o_addr[13] o_addr[14] _0319_ _0349_ _0256_ vssd1 vssd1 vccd1 vccd1 _0358_
+ sky130_fd_sc_hd__a41o_1
X_0773_ o_pc[5] _0253_ _0294_ o_pc_change _0297_ vssd1 vssd1 vccd1 vccd1 o_pc_next[5]
+ sky130_fd_sc_hd__a221o_4
X_1110_ clknet_4_6_0_i_clk u_buf.g_data\[0\].d_next\[17\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[0\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_1041_ clknet_4_5_0_i_clk u_buf.g_data\[2\].d_next\[14\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_0825_ o_pc[5] _0287_ _0324_ _0342_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__and4_1
X_0756_ o_addr[2] o_addr[3] o_addr[4] vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__a21o_1
X_0687_ u_buf.data\[1\]\[16\] _0222_ _0231_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[16\]
+ sky130_fd_sc_hd__a21o_1
X_0541_ u_buf.data\[3\]\[21\] _0143_ _0137_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__and3_1
X_0610_ u_buf.data\[1\]\[17\] _0178_ _0175_ i_instruction[17] _0185_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[1\].d_next\[17\] sky130_fd_sc_hd__a221o_1
X_0472_ u_buf.data\[0\]\[13\] u_buf.latch_hi\[13\] _0067_ vssd1 vssd1 vccd1 vccd1
+ _0100_ sky130_fd_sc_hd__mux2_1
X_1024_ clknet_4_12_0_i_clk u_buf.g_data\[3\].d_next\[30\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_0808_ o_addr[10] _0319_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__nand2_1
X_0739_ u_buf.data\[0\]\[0\] u_buf.data\[0\]\[1\] o_pc[1] vssd1 vssd1 vccd1 vccd1
+ _0267_ sky130_fd_sc_hd__a21o_1
X_0524_ u_buf.data\[2\]\[14\] _0127_ _0128_ i_instruction[14] _0134_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[14\] sky130_fd_sc_hd__a221o_1
X_0455_ _0091_ vssd1 vssd1 vccd1 vccd1 o_instruction[4] sky130_fd_sc_hd__buf_2
X_1007_ clknet_4_7_0_i_clk u_buf.g_data\[3\].d_next\[13\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_0438_ _0082_ vssd1 vssd1 vccd1 vccd1 o_instruction[28] sky130_fd_sc_hd__buf_2
X_0507_ u_buf.data\[2\]\[7\] _0109_ _0112_ i_instruction[7] _0124_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[7\] sky130_fd_sc_hd__a221o_1
X_0987_ _0060_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__clkbuf_1
X_0841_ o_pc[13] _0252_ _0354_ o_pc_change _0357_ vssd1 vssd1 vccd1 vccd1 o_pc_next[13]
+ sky130_fd_sc_hd__a221o_4
X_0772_ _0295_ _0296_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__nor2_1
X_0910_ _0387_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__clkbuf_1
X_1040_ clknet_4_7_0_i_clk u_buf.g_data\[2\].d_next\[13\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_0755_ o_pc[3] _0253_ _0278_ o_pc_change _0281_ vssd1 vssd1 vccd1 vccd1 o_pc_next[3]
+ sky130_fd_sc_hd__a221o_4
X_0824_ o_pc[9] o_pc[10] o_pc[11] o_pc[12] vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__and4_1
X_0686_ i_instruction[16] _0223_ _0224_ u_buf.data\[0\]\[16\] vssd1 vssd1 vccd1 vccd1
+ _0231_ sky130_fd_sc_hd__a22o_1
X_1169_ clknet_4_10_0_i_clk o_pc_next[13] vssd1 vssd1 vccd1 vccd1 o_pc[13] sky130_fd_sc_hd__dfxtp_4
X_0540_ u_buf.data\[2\]\[20\] _0141_ _0142_ i_instruction[20] _0144_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[20\] sky130_fd_sc_hd__a221o_1
X_0471_ _0099_ vssd1 vssd1 vccd1 vccd1 o_instruction[12] sky130_fd_sc_hd__buf_2
X_1023_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[29\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_0738_ _0068_ _0253_ _0260_ _0266_ vssd1 vssd1 vccd1 vccd1 o_pc_next[1] sky130_fd_sc_hd__a211o_4
X_0807_ o_pc[9] _0253_ _0323_ o_pc_change _0327_ vssd1 vssd1 vccd1 vccd1 o_pc_next[9]
+ sky130_fd_sc_hd__a221o_4
X_0669_ i_instruction[9] _0209_ _0211_ u_buf.data\[0\]\[9\] vssd1 vssd1 vccd1 vccd1
+ _0221_ sky130_fd_sc_hd__a22o_1
X_0523_ u_buf.data\[3\]\[14\] _0129_ _0123_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__and3_1
X_0454_ u_buf.data\[0\]\[4\] u_buf.latch_hi\[4\] _0088_ vssd1 vssd1 vccd1 vccd1 _0091_
+ sky130_fd_sc_hd__mux2_1
X_1006_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[12\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_0506_ u_buf.data\[3\]\[7\] _0113_ _0123_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__and3_1
X_0437_ u_buf.data\[0\]\[28\] u_buf.data\[0\]\[12\] _0077_ vssd1 vssd1 vccd1 vccd1
+ _0082_ sky130_fd_sc_hd__mux2_1
X_0986_ u_buf.data\[0\]\[30\] u_buf.latch_hi\[14\] _0250_ vssd1 vssd1 vccd1 vccd1
+ _0060_ sky130_fd_sc_hd__mux2_1
X_0840_ _0263_ _0355_ _0356_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__and3_1
X_0771_ o_pc[5] _0287_ _0264_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__o21ai_1
X_0969_ _0051_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__clkbuf_1
X_0754_ _0264_ _0279_ _0280_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__and3_1
X_0823_ o_pc[11] _0252_ _0338_ o_pc_change _0341_ vssd1 vssd1 vccd1 vccd1 o_pc_next[11]
+ sky130_fd_sc_hd__a221o_4
X_0685_ u_buf.data\[1\]\[15\] _0222_ _0230_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[15\]
+ sky130_fd_sc_hd__a21o_1
X_1168_ clknet_4_10_0_i_clk o_pc_next[12] vssd1 vssd1 vccd1 vccd1 o_pc[12] sky130_fd_sc_hd__dfxtp_4
X_1099_ clknet_4_0_0_i_clk u_buf.g_data\[0\].d_next\[6\] vssd1 vssd1 vccd1 vccd1 u_buf.data\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_0470_ u_buf.data\[0\]\[12\] u_buf.latch_hi\[12\] _0067_ vssd1 vssd1 vccd1 vccd1
+ _0099_ sky130_fd_sc_hd__mux2_1
X_1022_ clknet_4_15_0_i_clk u_buf.g_data\[3\].d_next\[28\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_0737_ _0067_ _0261_ _0264_ _0265_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__o211a_1
X_0806_ _0325_ _0263_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__and3b_1
X_0668_ u_buf.data\[1\]\[8\] _0208_ _0220_ vssd1 vssd1 vccd1 vccd1 u_buf.g_data\[0\].d_next\[8\]
+ sky130_fd_sc_hd__a21o_1
X_0599_ u_buf.data\[2\]\[12\] _0173_ _0176_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__and3_1
X_0522_ u_buf.data\[2\]\[13\] _0127_ _0128_ i_instruction[13] _0133_ vssd1 vssd1 vccd1
+ vccd1 u_buf.g_data\[2\].d_next\[13\] sky130_fd_sc_hd__a221o_1
X_0453_ _0090_ vssd1 vssd1 vccd1 vccd1 o_instruction[3] sky130_fd_sc_hd__buf_2
X_1005_ clknet_4_5_0_i_clk u_buf.g_data\[3\].d_next\[11\] vssd1 vssd1 vccd1 vccd1
+ u_buf.data\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_0505_ _0107_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__clkbuf_2
X_0436_ _0081_ vssd1 vssd1 vccd1 vccd1 o_instruction[27] sky130_fd_sc_hd__buf_2
.ends

