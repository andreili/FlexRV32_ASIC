* NGSPICE file created from rv_write.ext - technology: sky130A


X_363_ _165_ VSS VSS VCC VCC _029_ sky130_fd_sc_hd__clkbuf_1
X_294_ i_data[20] _118_ _127_ _054_ _055_ VSS VSS VCC VCC _128_ sky130_fd_sc_hd__a221o_1
X_346_ _156_ VSS VSS VCC VCC _021_ sky130_fd_sc_hd__clkbuf_1
X_415_ clknet_2_3__leaf_i_clk _027_ VSS VSS VCC VCC alu_result\[24\] sky130_fd_sc_hd__dfxtp_1
X_277_ i_data[9] i_data[25] _048_ VSS VSS VCC VCC _114_ sky130_fd_sc_hd__mux2_1
X_200_ _046_ _061_ _062_ _054_ VSS VSS VCC VCC _063_ sky130_fd_sc_hd__a22o_2
X_329_ _147_ VSS VSS VCC VCC _013_ sky130_fd_sc_hd__clkbuf_1
X_362_ i_alu_result[26] alu_result\[26\] _163_ VSS VSS VCC VCC _165_ sky130_fd_sc_hd__mux2_1
X_293_ i_data[12] i_data[28] _052_ VSS VSS VCC VCC _127_ sky130_fd_sc_hd__mux2_1
X_345_ i_alu_result[18] alu_result\[18\] _152_ VSS VSS VCC VCC _156_ sky130_fd_sc_hd__mux2_1
X_414_ clknet_2_3__leaf_i_clk _026_ VSS VSS VCC VCC alu_result\[23\] sky130_fd_sc_hd__dfxtp_1
X_276_ _043_ _111_ _113_ VSS VSS VCC VCC o_data[0] sky130_fd_sc_hd__a21o_2
X_259_ _098_ alu_result\[25\] _092_ _103_ VSS VSS VCC VCC o_data[25] sky130_fd_sc_hd__o22a_2
X_328_ i_alu_result[10] alu_result\[10\] _141_ VSS VSS VCC VCC _147_ sky130_fd_sc_hd__mux2_1
X_361_ _164_ VSS VSS VCC VCC _028_ sky130_fd_sc_hd__clkbuf_1
X_292_ i_data[4] _116_ VSS VSS VCC VCC _126_ sky130_fd_sc_hd__and2_1
X_344_ _155_ VSS VSS VCC VCC _020_ sky130_fd_sc_hd__clkbuf_1
X_413_ clknet_2_3__leaf_i_clk _025_ VSS VSS VCC VCC alu_result\[22\] sky130_fd_sc_hd__dfxtp_1
X_275_ _055_ alu_result\[0\] _054_ _112_ VSS VSS VCC VCC _113_ sky130_fd_sc_hd__a22o_1
X_258_ i_data[25] _093_ VSS VSS VCC VCC _103_ sky130_fd_sc_hd__and2_1
X_327_ _146_ VSS VSS VCC VCC _012_ sky130_fd_sc_hd__clkbuf_1
X_189_ i_data[14] i_data[30] _052_ VSS VSS VCC VCC _053_ sky130_fd_sc_hd__mux2_1
X_360_ i_alu_result[25] alu_result\[25\] _163_ VSS VSS VCC VCC _164_ sky130_fd_sc_hd__mux2_1
X_291_ _042_ alu_result\[3\] _123_ _125_ VSS VSS VCC VCC o_data[3] sky130_fd_sc_hd__o22a_2
X_412_ clknet_2_3__leaf_i_clk _024_ VSS VSS VCC VCC alu_result\[21\] sky130_fd_sc_hd__dfxtp_1
X_343_ i_alu_result[17] alu_result\[17\] _152_ VSS VSS VCC VCC _155_ sky130_fd_sc_hd__mux2_1
X_274_ i_data[8] i_data[24] _048_ VSS VSS VCC VCC _112_ sky130_fd_sc_hd__mux2_1
X_257_ _098_ alu_result\[24\] _092_ _102_ VSS VSS VCC VCC o_data[24] sky130_fd_sc_hd__o22a_2
X_326_ i_alu_result[9] alu_result\[9\] _141_ VSS VSS VCC VCC _146_ sky130_fd_sc_hd__mux2_1
X_188_ alu_result\[1\] VSS VSS VCC VCC _052_ sky130_fd_sc_hd__buf_2
X_309_ i_alu_result[1] _048_ _132_ VSS VSS VCC VCC _137_ sky130_fd_sc_hd__mux2_1
X_290_ i_data[19] _118_ _124_ _054_ _055_ VSS VSS VCC VCC _125_ sky130_fd_sc_hd__a221o_1
X_411_ clknet_2_2__leaf_i_clk _023_ VSS VSS VCC VCC alu_result\[20\] sky130_fd_sc_hd__dfxtp_1
X_342_ _154_ VSS VSS VCC VCC _019_ sky130_fd_sc_hd__clkbuf_1
X_273_ i_data[0] _051_ _110_ _047_ VSS VSS VCC VCC _111_ sky130_fd_sc_hd__a22o_1
X_187_ _050_ VSS VSS VCC VCC _051_ sky130_fd_sc_hd__clkbuf_2
X_325_ _145_ VSS VSS VCC VCC _011_ sky130_fd_sc_hd__clkbuf_1
X_256_ i_data[24] _093_ VSS VSS VCC VCC _102_ sky130_fd_sc_hd__and2_1
X_308_ _136_ VSS VSS VCC VCC _003_ sky130_fd_sc_hd__clkbuf_1
X_239_ _043_ alu_result\[16\] _089_ _092_ VSS VSS VCC VCC o_data[16] sky130_fd_sc_hd__o22a_2
Xclkbuf_0_i_clk i_clk VSS VSS VCC VCC clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_410_ clknet_2_3__leaf_i_clk _022_ VSS VSS VCC VCC alu_result\[19\] sky130_fd_sc_hd__dfxtp_1
X_341_ i_alu_result[16] alu_result\[16\] _152_ VSS VSS VCC VCC _154_ sky130_fd_sc_hd__mux2_1
X_272_ i_data[0] i_data[16] _048_ VSS VSS VCC VCC _110_ sky130_fd_sc_hd__mux2_1
X_186_ funct3\[0\] funct3\[2\] funct3\[1\] VSS VSS VCC VCC _050_ sky130_fd_sc_hd__nor3b_1
X_324_ i_alu_result[8] alu_result\[8\] _141_ VSS VSS VCC VCC _145_ sky130_fd_sc_hd__mux2_1
X_255_ _098_ alu_result\[23\] _092_ _101_ VSS VSS VCC VCC o_data[23] sky130_fd_sc_hd__o22a_2
X_307_ i_alu_result[0] alu_result\[0\] _132_ VSS VSS VCC VCC _136_ sky130_fd_sc_hd__mux2_1
X_238_ _091_ VSS VSS VCC VCC _092_ sky130_fd_sc_hd__buf_2
X_340_ _153_ VSS VSS VCC VCC _018_ sky130_fd_sc_hd__clkbuf_1
X_271_ _042_ alu_result\[31\] _091_ _109_ VSS VSS VCC VCC o_data[31] sky130_fd_sc_hd__o22a_2
X_254_ i_data[23] _093_ VSS VSS VCC VCC _101_ sky130_fd_sc_hd__and2_1
X_323_ _144_ VSS VSS VCC VCC _010_ sky130_fd_sc_hd__clkbuf_1
X_185_ i_data[6] i_data[22] _048_ VSS VSS VCC VCC _049_ sky130_fd_sc_hd__mux2_1
X_306_ _135_ VSS VSS VCC VCC _002_ sky130_fd_sc_hd__clkbuf_1
X_237_ _065_ _063_ _090_ VSS VSS VCC VCC _091_ sky130_fd_sc_hd__a21o_1
X_270_ i_data[31] _051_ VSS VSS VCC VCC _109_ sky130_fd_sc_hd__and2_1
X_399_ clknet_2_0__leaf_i_clk _011_ VSS VSS VCC VCC alu_result\[8\] sky130_fd_sc_hd__dfxtp_1
X_322_ i_alu_result[7] alu_result\[7\] _141_ VSS VSS VCC VCC _144_ sky130_fd_sc_hd__mux2_1
X_184_ alu_result\[1\] VSS VSS VCC VCC _048_ sky130_fd_sc_hd__clkbuf_4
X_253_ _098_ alu_result\[22\] _092_ _100_ VSS VSS VCC VCC o_data[22] sky130_fd_sc_hd__o22a_2
X_305_ i_funct3[2] funct3\[2\] _132_ VSS VSS VCC VCC _135_ sky130_fd_sc_hd__mux2_1
X_236_ _065_ _045_ _062_ _055_ VSS VSS VCC VCC _090_ sky130_fd_sc_hd__a31o_1
X_219_ _077_ VSS VSS VCC VCC o_data[11] sky130_fd_sc_hd__buf_2
X_398_ clknet_2_0__leaf_i_clk _010_ VSS VSS VCC VCC alu_result\[7\] sky130_fd_sc_hd__dfxtp_1
X_252_ i_data[22] _093_ VSS VSS VCC VCC _100_ sky130_fd_sc_hd__and2_1
X_183_ _045_ _046_ VSS VSS VCC VCC _047_ sky130_fd_sc_hd__or2_1
X_321_ _143_ VSS VSS VCC VCC _009_ sky130_fd_sc_hd__clkbuf_1
X_304_ _134_ VSS VSS VCC VCC _001_ sky130_fd_sc_hd__clkbuf_1
X_235_ i_data[16] _051_ VSS VSS VCC VCC _089_ sky130_fd_sc_hd__and2_1
X_218_ alu_result\[11\] _076_ res_src\[2\] VSS VSS VCC VCC _077_ sky130_fd_sc_hd__mux2_1
X_397_ clknet_2_0__leaf_i_clk _009_ VSS VSS VCC VCC alu_result\[6\] sky130_fd_sc_hd__dfxtp_1
X_182_ funct3\[1\] funct3\[0\] alu_result\[0\] VSS VSS VCC VCC _046_ sky130_fd_sc_hd__nor3_1
X_251_ _098_ alu_result\[21\] _092_ _099_ VSS VSS VCC VCC o_data[21] sky130_fd_sc_hd__o22a_2
X_320_ i_alu_result[6] alu_result\[6\] _141_ VSS VSS VCC VCC _143_ sky130_fd_sc_hd__mux2_1
X_303_ i_funct3[1] funct3\[1\] _132_ VSS VSS VCC VCC _134_ sky130_fd_sc_hd__mux2_1
X_234_ _043_ alu_result\[15\] _088_ VSS VSS VCC VCC o_data[15] sky130_fd_sc_hd__o21a_2
Xclkbuf_2_2__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_2__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_217_ _065_ _063_ _059_ i_data[11] _075_ VSS VSS VCC VCC _076_ sky130_fd_sc_hd__a221o_1
X_396_ clknet_2_1__leaf_i_clk _008_ VSS VSS VCC VCC alu_result\[5\] sky130_fd_sc_hd__dfxtp_1
X_181_ _044_ VSS VSS VCC VCC _045_ sky130_fd_sc_hd__buf_2
X_250_ i_data[21] _093_ VSS VSS VCC VCC _099_ sky130_fd_sc_hd__and2_1
X_379_ _173_ VSS VSS VCC VCC _037_ sky130_fd_sc_hd__clkbuf_1
X_302_ _133_ VSS VSS VCC VCC _000_ sky130_fd_sc_hd__clkbuf_1
X_233_ _065_ _063_ _087_ VSS VSS VCC VCC _088_ sky130_fd_sc_hd__a21o_1
X_216_ _052_ i_data[27] _045_ VSS VSS VCC VCC _075_ sky130_fd_sc_hd__and3_1
X_395_ clknet_2_0__leaf_i_clk _007_ VSS VSS VCC VCC alu_result\[4\] sky130_fd_sc_hd__dfxtp_1
X_180_ funct3\[1\] funct3\[0\] VSS VSS VCC VCC _044_ sky130_fd_sc_hd__and2b_1
X_378_ i_rd[0] o_rd[0] _163_ VSS VSS VCC VCC _173_ sky130_fd_sc_hd__mux2_1
X_301_ i_funct3[0] funct3\[0\] _132_ VSS VSS VCC VCC _133_ sky130_fd_sc_hd__mux2_1
X_232_ i_data[15] _051_ _062_ _045_ _055_ VSS VSS VCC VCC _087_ sky130_fd_sc_hd__a221o_1
X_215_ _074_ VSS VSS VCC VCC o_data[10] sky130_fd_sc_hd__buf_2
X_394_ clknet_2_0__leaf_i_clk _006_ VSS VSS VCC VCC alu_result\[3\] sky130_fd_sc_hd__dfxtp_1
X_377_ _172_ VSS VSS VCC VCC _036_ sky130_fd_sc_hd__clkbuf_1
X_300_ i_flush VSS VSS VCC VCC _132_ sky130_fd_sc_hd__clkbuf_4
X_231_ _086_ VSS VSS VCC VCC o_data[14] sky130_fd_sc_hd__buf_2
X_429_ clknet_2_3__leaf_i_clk _041_ VSS VSS VCC VCC o_rd[4] sky130_fd_sc_hd__dfxtp_2
X_214_ alu_result\[10\] _073_ _042_ VSS VSS VCC VCC _074_ sky130_fd_sc_hd__mux2_1
X_393_ clknet_2_1__leaf_i_clk _005_ VSS VSS VCC VCC alu_result\[2\] sky130_fd_sc_hd__dfxtp_1
X_376_ _132_ i_reg_write VSS VSS VCC VCC _172_ sky130_fd_sc_hd__and2b_1
X_230_ alu_result\[14\] _085_ res_src\[2\] VSS VSS VCC VCC _086_ sky130_fd_sc_hd__mux2_1
X_359_ i_flush VSS VSS VCC VCC _163_ sky130_fd_sc_hd__clkbuf_4
X_428_ clknet_2_3__leaf_i_clk _040_ VSS VSS VCC VCC o_rd[3] sky130_fd_sc_hd__dfxtp_2
X_213_ _065_ _063_ _059_ i_data[10] _072_ VSS VSS VCC VCC _073_ sky130_fd_sc_hd__a221o_1
X_392_ clknet_2_1__leaf_i_clk _004_ VSS VSS VCC VCC alu_result\[1\] sky130_fd_sc_hd__dfxtp_1
X_375_ _171_ VSS VSS VCC VCC _035_ sky130_fd_sc_hd__clkbuf_1
X_358_ _162_ VSS VSS VCC VCC _027_ sky130_fd_sc_hd__clkbuf_1
X_427_ clknet_2_1__leaf_i_clk _039_ VSS VSS VCC VCC o_rd[2] sky130_fd_sc_hd__dfxtp_2
X_289_ i_data[11] i_data[27] _048_ VSS VSS VCC VCC _124_ sky130_fd_sc_hd__mux2_1
X_212_ _052_ i_data[26] _045_ VSS VSS VCC VCC _072_ sky130_fd_sc_hd__and3_1
X_391_ clknet_2_2__leaf_i_clk _003_ VSS VSS VCC VCC alu_result\[0\] sky130_fd_sc_hd__dfxtp_1
X_374_ _132_ i_res_src[2] VSS VSS VCC VCC _171_ sky130_fd_sc_hd__and2b_1
X_357_ i_alu_result[24] alu_result\[24\] _152_ VSS VSS VCC VCC _162_ sky130_fd_sc_hd__mux2_1
X_426_ clknet_2_3__leaf_i_clk _038_ VSS VSS VCC VCC o_rd[1] sky130_fd_sc_hd__dfxtp_2
X_288_ i_data[3] _116_ VSS VSS VCC VCC _123_ sky130_fd_sc_hd__and2_1
X_211_ _071_ VSS VSS VCC VCC o_data[9] sky130_fd_sc_hd__buf_2
X_409_ clknet_2_3__leaf_i_clk _021_ VSS VSS VCC VCC alu_result\[18\] sky130_fd_sc_hd__dfxtp_1
X_390_ clknet_2_0__leaf_i_clk _002_ VSS VSS VCC VCC funct3\[2\] sky130_fd_sc_hd__dfxtp_1
X_373_ _170_ VSS VSS VCC VCC _034_ sky130_fd_sc_hd__clkbuf_1
X_356_ _161_ VSS VSS VCC VCC _026_ sky130_fd_sc_hd__clkbuf_1
X_425_ clknet_2_1__leaf_i_clk _037_ VSS VSS VCC VCC o_rd[0] sky130_fd_sc_hd__dfxtp_2
X_287_ _042_ alu_result\[2\] _120_ _122_ VSS VSS VCC VCC o_data[2] sky130_fd_sc_hd__o22a_2
X_408_ clknet_2_3__leaf_i_clk _020_ VSS VSS VCC VCC alu_result\[17\] sky130_fd_sc_hd__dfxtp_1
X_210_ alu_result\[9\] _070_ _042_ VSS VSS VCC VCC _071_ sky130_fd_sc_hd__mux2_1
X_339_ i_alu_result[15] alu_result\[15\] _152_ VSS VSS VCC VCC _153_ sky130_fd_sc_hd__mux2_1
X_372_ i_alu_result[31] alu_result\[31\] _163_ VSS VSS VCC VCC _170_ sky130_fd_sc_hd__mux2_1
X_355_ i_alu_result[23] alu_result\[23\] _152_ VSS VSS VCC VCC _161_ sky130_fd_sc_hd__mux2_1
X_424_ clknet_2_0__leaf_i_clk _036_ VSS VSS VCC VCC o_write_op sky130_fd_sc_hd__dfxtp_2
X_286_ i_data[18] _118_ _121_ _054_ _055_ VSS VSS VCC VCC _122_ sky130_fd_sc_hd__a221o_1
X_338_ i_flush VSS VSS VCC VCC _152_ sky130_fd_sc_hd__clkbuf_4
X_407_ clknet_2_2__leaf_i_clk _019_ VSS VSS VCC VCC alu_result\[16\] sky130_fd_sc_hd__dfxtp_1
X_269_ _098_ alu_result\[30\] _091_ _108_ VSS VSS VCC VCC o_data[30] sky130_fd_sc_hd__o22a_2
X_371_ _169_ VSS VSS VCC VCC _033_ sky130_fd_sc_hd__clkbuf_1
X_354_ _160_ VSS VSS VCC VCC _025_ sky130_fd_sc_hd__clkbuf_1
X_423_ clknet_2_1__leaf_i_clk _035_ VSS VSS VCC VCC res_src\[2\] sky130_fd_sc_hd__dfxtp_2
X_285_ i_data[10] i_data[26] _048_ VSS VSS VCC VCC _121_ sky130_fd_sc_hd__mux2_1
X_406_ clknet_2_2__leaf_i_clk _018_ VSS VSS VCC VCC alu_result\[15\] sky130_fd_sc_hd__dfxtp_1
X_337_ _151_ VSS VSS VCC VCC _017_ sky130_fd_sc_hd__clkbuf_1
X_268_ i_data[30] _051_ VSS VSS VCC VCC _108_ sky130_fd_sc_hd__and2_1
X_199_ i_data[15] i_data[31] alu_result\[1\] VSS VSS VCC VCC _062_ sky130_fd_sc_hd__mux2_1
X_370_ i_alu_result[30] alu_result\[30\] _163_ VSS VSS VCC VCC _169_ sky130_fd_sc_hd__mux2_1
X_353_ i_alu_result[22] alu_result\[22\] _152_ VSS VSS VCC VCC _160_ sky130_fd_sc_hd__mux2_1
X_422_ clknet_2_1__leaf_i_clk _034_ VSS VSS VCC VCC alu_result\[31\] sky130_fd_sc_hd__dfxtp_1
X_284_ i_data[2] _116_ VSS VSS VCC VCC _120_ sky130_fd_sc_hd__and2_1
X_405_ clknet_2_2__leaf_i_clk _017_ VSS VSS VCC VCC alu_result\[14\] sky130_fd_sc_hd__dfxtp_1
X_336_ i_alu_result[14] alu_result\[14\] _141_ VSS VSS VCC VCC _151_ sky130_fd_sc_hd__mux2_1
X_267_ _098_ alu_result\[29\] _091_ _107_ VSS VSS VCC VCC o_data[29] sky130_fd_sc_hd__o22a_2
X_198_ i_data[7] i_data[23] alu_result\[1\] VSS VSS VCC VCC _061_ sky130_fd_sc_hd__mux2_1
X_319_ _142_ VSS VSS VCC VCC _008_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_1__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_1__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_421_ clknet_2_1__leaf_i_clk _033_ VSS VSS VCC VCC alu_result\[30\] sky130_fd_sc_hd__dfxtp_1
X_352_ _159_ VSS VSS VCC VCC _024_ sky130_fd_sc_hd__clkbuf_1
X_283_ _043_ _117_ _119_ VSS VSS VCC VCC o_data[1] sky130_fd_sc_hd__a21o_2
X_335_ _150_ VSS VSS VCC VCC _016_ sky130_fd_sc_hd__clkbuf_1
X_404_ clknet_2_2__leaf_i_clk _016_ VSS VSS VCC VCC alu_result\[13\] sky130_fd_sc_hd__dfxtp_1
X_266_ i_data[29] _051_ VSS VSS VCC VCC _107_ sky130_fd_sc_hd__and2_1
X_197_ _048_ i_data[23] _045_ _055_ VSS VSS VCC VCC _060_ sky130_fd_sc_hd__a31o_1
X_249_ _042_ VSS VSS VCC VCC _098_ sky130_fd_sc_hd__buf_2
X_318_ i_alu_result[5] alu_result\[5\] _141_ VSS VSS VCC VCC _142_ sky130_fd_sc_hd__mux2_1
X_351_ i_alu_result[21] alu_result\[21\] _152_ VSS VSS VCC VCC _159_ sky130_fd_sc_hd__mux2_1
X_420_ clknet_2_1__leaf_i_clk _032_ VSS VSS VCC VCC alu_result\[29\] sky130_fd_sc_hd__dfxtp_1
X_282_ _048_ _055_ i_data[17] _118_ VSS VSS VCC VCC _119_ sky130_fd_sc_hd__a22o_1
X_334_ i_alu_result[13] alu_result\[13\] _141_ VSS VSS VCC VCC _150_ sky130_fd_sc_hd__mux2_1
X_403_ clknet_2_2__leaf_i_clk _015_ VSS VSS VCC VCC alu_result\[12\] sky130_fd_sc_hd__dfxtp_1
X_196_ _050_ _058_ VSS VSS VCC VCC _059_ sky130_fd_sc_hd__nand2b_2
X_265_ _098_ alu_result\[28\] _091_ _106_ VSS VSS VCC VCC o_data[28] sky130_fd_sc_hd__o22a_2
X_317_ i_flush VSS VSS VCC VCC _141_ sky130_fd_sc_hd__clkbuf_4
X_179_ _042_ VSS VSS VCC VCC _043_ sky130_fd_sc_hd__buf_2
X_248_ _043_ alu_result\[20\] _092_ _097_ VSS VSS VCC VCC o_data[20] sky130_fd_sc_hd__o22a_2
X_350_ _158_ VSS VSS VCC VCC _023_ sky130_fd_sc_hd__clkbuf_1
X_281_ _045_ _046_ _048_ VSS VSS VCC VCC _118_ sky130_fd_sc_hd__o21a_1
X_333_ _149_ VSS VSS VCC VCC _015_ sky130_fd_sc_hd__clkbuf_1
X_402_ clknet_2_2__leaf_i_clk _014_ VSS VSS VCC VCC alu_result\[11\] sky130_fd_sc_hd__dfxtp_1
X_195_ alu_result\[1\] funct3\[1\] funct3\[0\] VSS VSS VCC VCC _058_ sky130_fd_sc_hd__or3b_1
X_264_ i_data[28] _051_ VSS VSS VCC VCC _106_ sky130_fd_sc_hd__and2_1
X_316_ _140_ VSS VSS VCC VCC _007_ sky130_fd_sc_hd__clkbuf_1
X_247_ i_data[20] _093_ VSS VSS VCC VCC _097_ sky130_fd_sc_hd__and2_1
X_178_ res_src\[2\] VSS VSS VCC VCC _042_ sky130_fd_sc_hd__buf_2
X_280_ _054_ _114_ _116_ i_data[1] VSS VSS VCC VCC _117_ sky130_fd_sc_hd__a22o_1
X_332_ i_alu_result[12] alu_result\[12\] _141_ VSS VSS VCC VCC _149_ sky130_fd_sc_hd__mux2_1
X_401_ clknet_2_1__leaf_i_clk _013_ VSS VSS VCC VCC alu_result\[10\] sky130_fd_sc_hd__dfxtp_1
X_263_ _098_ alu_result\[27\] _091_ _105_ VSS VSS VCC VCC o_data[27] sky130_fd_sc_hd__o22a_2
X_194_ alu_result\[6\] _043_ _057_ VSS VSS VCC VCC o_data[6] sky130_fd_sc_hd__o21a_2
X_315_ i_alu_result[4] alu_result\[4\] _132_ VSS VSS VCC VCC _140_ sky130_fd_sc_hd__mux2_1
X_246_ _043_ alu_result\[19\] _092_ _096_ VSS VSS VCC VCC o_data[19] sky130_fd_sc_hd__o22a_2
X_229_ _065_ _063_ _059_ i_data[14] _084_ VSS VSS VCC VCC _085_ sky130_fd_sc_hd__a221o_1
X_331_ _148_ VSS VSS VCC VCC _014_ sky130_fd_sc_hd__clkbuf_1
X_400_ clknet_2_0__leaf_i_clk _012_ VSS VSS VCC VCC alu_result\[9\] sky130_fd_sc_hd__dfxtp_1
X_262_ i_data[27] _051_ VSS VSS VCC VCC _105_ sky130_fd_sc_hd__and2_1
X_193_ _047_ _049_ _056_ VSS VSS VCC VCC _057_ sky130_fd_sc_hd__a21o_1
X_314_ _139_ VSS VSS VCC VCC _006_ sky130_fd_sc_hd__clkbuf_1
X_245_ i_data[19] _093_ VSS VSS VCC VCC _096_ sky130_fd_sc_hd__and2_1
X_228_ _052_ i_data[30] _044_ VSS VSS VCC VCC _084_ sky130_fd_sc_hd__and3_1
X_330_ i_alu_result[11] alu_result\[11\] _141_ VSS VSS VCC VCC _148_ sky130_fd_sc_hd__mux2_1
X_261_ _098_ alu_result\[26\] _091_ _104_ VSS VSS VCC VCC o_data[26] sky130_fd_sc_hd__o22a_2
X_192_ i_data[6] _051_ _053_ _054_ _055_ VSS VSS VCC VCC _056_ sky130_fd_sc_hd__a221o_1
X_313_ i_alu_result[3] alu_result\[3\] _132_ VSS VSS VCC VCC _139_ sky130_fd_sc_hd__mux2_1
X_244_ _043_ alu_result\[18\] _092_ _095_ VSS VSS VCC VCC o_data[18] sky130_fd_sc_hd__o22a_2
X_227_ _083_ VSS VSS VCC VCC o_data[13] sky130_fd_sc_hd__buf_2
X_260_ i_data[26] _093_ VSS VSS VCC VCC _104_ sky130_fd_sc_hd__and2_1
X_389_ clknet_2_0__leaf_i_clk _001_ VSS VSS VCC VCC funct3\[1\] sky130_fd_sc_hd__dfxtp_2
X_191_ res_src\[2\] VSS VSS VCC VCC _055_ sky130_fd_sc_hd__inv_2
X_312_ _138_ VSS VSS VCC VCC _005_ sky130_fd_sc_hd__clkbuf_1
X_243_ i_data[18] _093_ VSS VSS VCC VCC _095_ sky130_fd_sc_hd__and2_1
X_226_ alu_result\[13\] _082_ res_src\[2\] VSS VSS VCC VCC _083_ sky130_fd_sc_hd__mux2_1
X_209_ _065_ _063_ _059_ i_data[9] _069_ VSS VSS VCC VCC _070_ sky130_fd_sc_hd__a221o_1
X_190_ funct3\[1\] funct3\[0\] alu_result\[0\] VSS VSS VCC VCC _054_ sky130_fd_sc_hd__nor3b_4
X_388_ clknet_2_0__leaf_i_clk _000_ VSS VSS VCC VCC funct3\[0\] sky130_fd_sc_hd__dfxtp_2
X_311_ i_alu_result[2] alu_result\[2\] _132_ VSS VSS VCC VCC _138_ sky130_fd_sc_hd__mux2_1
X_242_ _043_ alu_result\[17\] _092_ _094_ VSS VSS VCC VCC o_data[17] sky130_fd_sc_hd__o22a_2
X_225_ _065_ _063_ _059_ i_data[13] _081_ VSS VSS VCC VCC _082_ sky130_fd_sc_hd__a221o_1
X_208_ _052_ i_data[25] _045_ VSS VSS VCC VCC _069_ sky130_fd_sc_hd__and3_1
X_387_ _177_ VSS VSS VCC VCC _041_ sky130_fd_sc_hd__clkbuf_1
X_310_ _137_ VSS VSS VCC VCC _004_ sky130_fd_sc_hd__clkbuf_1
X_241_ i_data[17] _093_ VSS VSS VCC VCC _094_ sky130_fd_sc_hd__and2_1
X_224_ _052_ i_data[29] _044_ VSS VSS VCC VCC _081_ sky130_fd_sc_hd__and3_1
X_207_ _068_ VSS VSS VCC VCC o_data[8] sky130_fd_sc_hd__buf_2
X_386_ i_rd[4] o_rd[4] i_flush VSS VSS VCC VCC _177_ sky130_fd_sc_hd__mux2_1
X_240_ _051_ VSS VSS VCC VCC _093_ sky130_fd_sc_hd__clkbuf_2
X_369_ _168_ VSS VSS VCC VCC _032_ sky130_fd_sc_hd__clkbuf_1
X_223_ _080_ VSS VSS VCC VCC o_data[12] sky130_fd_sc_hd__buf_2
X_206_ alu_result\[8\] _067_ _042_ VSS VSS VCC VCC _068_ sky130_fd_sc_hd__mux2_1
X_385_ _176_ VSS VSS VCC VCC _040_ sky130_fd_sc_hd__clkbuf_1
X_368_ i_alu_result[29] alu_result\[29\] _163_ VSS VSS VCC VCC _168_ sky130_fd_sc_hd__mux2_1
X_299_ _042_ alu_result\[5\] _129_ _131_ VSS VSS VCC VCC o_data[5] sky130_fd_sc_hd__o22a_2
Xclkbuf_2_0__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_0__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_222_ alu_result\[12\] _079_ res_src\[2\] VSS VSS VCC VCC _080_ sky130_fd_sc_hd__mux2_1
X_205_ _065_ _063_ _059_ i_data[8] _066_ VSS VSS VCC VCC _067_ sky130_fd_sc_hd__a221o_1
X_384_ i_rd[3] o_rd[3] i_flush VSS VSS VCC VCC _176_ sky130_fd_sc_hd__mux2_1
X_367_ _167_ VSS VSS VCC VCC _031_ sky130_fd_sc_hd__clkbuf_1
X_298_ i_data[21] _118_ _130_ _054_ _055_ VSS VSS VCC VCC _131_ sky130_fd_sc_hd__a221o_1
X_221_ _065_ _063_ _059_ i_data[12] _078_ VSS VSS VCC VCC _079_ sky130_fd_sc_hd__a221o_1
X_419_ clknet_2_3__leaf_i_clk _031_ VSS VSS VCC VCC alu_result\[28\] sky130_fd_sc_hd__dfxtp_1
X_204_ _052_ i_data[24] _045_ VSS VSS VCC VCC _066_ sky130_fd_sc_hd__and3_1
X_383_ _175_ VSS VSS VCC VCC _039_ sky130_fd_sc_hd__clkbuf_1
X_366_ i_alu_result[28] alu_result\[28\] _163_ VSS VSS VCC VCC _167_ sky130_fd_sc_hd__mux2_1
X_297_ i_data[13] i_data[29] _052_ VSS VSS VCC VCC _130_ sky130_fd_sc_hd__mux2_1
X_220_ _052_ i_data[28] _045_ VSS VSS VCC VCC _078_ sky130_fd_sc_hd__and3_1
X_349_ i_alu_result[20] alu_result\[20\] _152_ VSS VSS VCC VCC _158_ sky130_fd_sc_hd__mux2_1
X_418_ clknet_2_1__leaf_i_clk _030_ VSS VSS VCC VCC alu_result\[27\] sky130_fd_sc_hd__dfxtp_1
X_203_ funct3\[2\] VSS VSS VCC VCC _065_ sky130_fd_sc_hd__inv_2
X_382_ i_rd[2] o_rd[2] _163_ VSS VSS VCC VCC _175_ sky130_fd_sc_hd__mux2_1
X_365_ _166_ VSS VSS VCC VCC _030_ sky130_fd_sc_hd__clkbuf_1
X_296_ i_data[5] _116_ VSS VSS VCC VCC _129_ sky130_fd_sc_hd__and2_1
X_348_ _157_ VSS VSS VCC VCC _022_ sky130_fd_sc_hd__clkbuf_1
X_417_ clknet_2_1__leaf_i_clk _029_ VSS VSS VCC VCC alu_result\[26\] sky130_fd_sc_hd__dfxtp_1
X_279_ _050_ _058_ _115_ VSS VSS VCC VCC _116_ sky130_fd_sc_hd__nand3b_2
X_202_ _043_ alu_result\[7\] _064_ VSS VSS VCC VCC o_data[7] sky130_fd_sc_hd__o21a_2
Xclkbuf_2_3__f_i_clk clknet_0_i_clk VSS VSS VCC VCC clknet_2_3__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_381_ _174_ VSS VSS VCC VCC _038_ sky130_fd_sc_hd__clkbuf_1
X_364_ i_alu_result[27] alu_result\[27\] _163_ VSS VSS VCC VCC _166_ sky130_fd_sc_hd__mux2_1
X_295_ _042_ alu_result\[4\] _126_ _128_ VSS VSS VCC VCC o_data[4] sky130_fd_sc_hd__o22a_2
X_347_ i_alu_result[19] alu_result\[19\] _152_ VSS VSS VCC VCC _157_ sky130_fd_sc_hd__mux2_1
X_416_ clknet_2_1__leaf_i_clk _028_ VSS VSS VCC VCC alu_result\[25\] sky130_fd_sc_hd__dfxtp_1
X_278_ alu_result\[1\] funct3\[1\] funct3\[0\] alu_result\[0\] VSS VSS VCC VCC
+ _115_ sky130_fd_sc_hd__or4_1
X_201_ i_data[7] _059_ _060_ _063_ VSS VSS VCC VCC _064_ sky130_fd_sc_hd__a211o_1
X_380_ i_rd[1] o_rd[1] _163_ VSS VSS VCC VCC _174_ sky130_fd_sc_hd__mux2_1
