* NGSPICE file created from rv_decode.ext - technology: sky130A

.subckt rv_decode
+ i_clk i_flush
+ i_instruction[0] i_instruction[1] i_instruction[2] i_instruction[3] i_instruction[4] i_instruction[5] i_instruction[6] i_instruction[7] i_instruction[8] i_instruction[9] i_instruction[10] i_instruction[11] i_instruction[12] i_instruction[13] i_instruction[14] i_instruction[15] i_instruction[16] i_instruction[17] i_instruction[18] i_instruction[19] i_instruction[20] i_instruction[21] i_instruction[22] i_instruction[23] i_instruction[24] i_instruction[25] i_instruction[26] i_instruction[27] i_instruction[28] i_instruction[29] i_instruction[30] i_instruction[31] 
+ i_pc[1] i_pc[2] i_pc[3] i_pc[4] i_pc[5] i_pc[6] i_pc[7] i_pc[8] i_pc[9] i_pc[10] i_pc[11] i_pc[12] i_pc[13] i_pc[14] i_pc[15] 
+ i_pc_next[1] i_pc_next[2] i_pc_next[3] i_pc_next[4] i_pc_next[5] i_pc_next[6] i_pc_next[7] i_pc_next[8] i_pc_next[9] i_pc_next[10] i_pc_next[11] i_pc_next[12] i_pc_next[13] i_pc_next[14] i_pc_next[15] 
+ i_ready i_stall
+ o_csr_idx[0] o_csr_idx[1] o_csr_idx[2] o_csr_idx[3] o_csr_idx[4] o_csr_idx[5] o_csr_idx[6] o_csr_idx[7] o_csr_idx[8] o_csr_idx[9] o_csr_idx[10] o_csr_idx[11] 
+ o_csr_imm[0] o_csr_imm[1] o_csr_imm[2] o_csr_imm[3] o_csr_imm[4] 
+ o_csr_pc_next[1] o_csr_pc_next[2] o_csr_pc_next[3] o_csr_pc_next[4] o_csr_pc_next[5] o_csr_pc_next[6] o_csr_pc_next[7] o_csr_pc_next[8] o_csr_pc_next[9] o_csr_pc_next[10] o_csr_pc_next[11] o_csr_pc_next[12] o_csr_pc_next[13] o_csr_pc_next[14] o_csr_pc_next[15] 
+ o_csr_clear o_csr_ebreak o_csr_read o_csr_set o_csr_write o_csr_imm_sel
+ o_imm_i[0] o_imm_i[1] o_imm_i[2] o_imm_i[3] o_imm_i[4] o_imm_i[5] o_imm_i[6] o_imm_i[7] o_imm_i[8] o_imm_i[9] o_imm_i[10] o_imm_i[11] o_imm_i[12] o_imm_i[13] o_imm_i[14] o_imm_i[15] o_imm_i[16] o_imm_i[17] o_imm_i[18] o_imm_i[19] o_imm_i[20] o_imm_i[21] o_imm_i[22] o_imm_i[23] o_imm_i[24] o_imm_i[25] o_imm_i[26] o_imm_i[27] o_imm_i[28] o_imm_i[29] o_imm_i[30] o_imm_i[31] 
+ o_alu_ctrl[0] o_alu_ctrl[1] o_alu_ctrl[2] o_alu_ctrl[3] o_alu_ctrl[4] 
+ o_funct3[0] o_funct3[1] o_funct3[2]
+ o_reg_write o_op1_src o_op2_src o_inst_branch o_inst_csr_req o_inst_jal o_inst_jalr o_inst_mret o_inst_store o_inst_supported
+ o_pc[1] o_pc[2] o_pc[3] o_pc[4] o_pc[5] o_pc[6] o_pc[7] o_pc[8] o_pc[9] o_pc[10] o_pc[11] o_pc[12] o_pc[13] o_pc[14] o_pc[15] 
+ o_pc_next[1] o_pc_next[2] o_pc_next[3] o_pc_next[4] o_pc_next[5] o_pc_next[6] o_pc_next[7] o_pc_next[8] o_pc_next[9] o_pc_next[10] o_pc_next[11] o_pc_next[12] o_pc_next[13] o_pc_next[14] o_pc_next[15] 
+ o_rd[0] o_rd[1] o_rd[2] o_rd[3] o_rd[4] 
+ o_rs1[0] o_rs1[1] o_rs1[2] o_rs1[3] o_rs1[4] 
+ o_rs2[0] o_rs2[1] o_rs2[2] o_rs2[3] o_rs2[4] 
+ o_res_src[0] o_res_src[1] o_res_src[2] 
+ vccd1 vssd1
X_0985_ clknet_3_4__leaf_i_clk _0014_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[15] sky130_fd_sc_hd__dfxtp_2
X_0770_ i_instruction[10] _0283_ _0292_ _0228_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__a211o_1
X_0968_ _0455_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__clkbuf_1
X_0899_ _0168_ _0403_ _0405_ _0406_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__or4_2
X_0822_ _0330_ _0338_ _0174_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__a21o_1
X_0753_ i_instruction[3] _0273_ _0277_ i_instruction[8] _0260_ vssd1 vssd1 vccd1 vccd1
+ _0278_ sky130_fd_sc_hd__a221o_1
X_0684_ _0214_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__buf_6
X_1021_ clknet_3_2__leaf_i_clk _0050_ vssd1 vssd1 vccd1 vccd1 o_pc[3] sky130_fd_sc_hd__dfxtp_2
X_0805_ _0172_ i_instruction[5] _0213_ _0322_ _0249_ vssd1 vssd1 vccd1 vccd1 _0323_
+ sky130_fd_sc_hd__a32o_1
X_0736_ i_instruction[12] _0223_ _0236_ _0249_ _0257_ vssd1 vssd1 vccd1 vccd1 _0262_
+ sky130_fd_sc_hd__a221o_1
X_0667_ _0170_ i_instruction[4] vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__nand2_4
X_0598_ _0146_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__buf_12
X_0521_ o_csr_idx[4] vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__inv_2
X_1004_ clknet_3_3__leaf_i_clk _0033_ vssd1 vssd1 vccd1 vccd1 o_csr_imm[2] sky130_fd_sc_hd__dfxtp_4
X_0719_ _0229_ _0245_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__nor2_1
X_0504_ instruction\[5\] _0075_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__nand2_1
X_0984_ clknet_3_7__leaf_i_clk _0013_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[14] sky130_fd_sc_hd__dfxtp_2
X_0967_ o_pc[14] i_pc[14] _0446_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__mux2_1
X_0898_ _0177_ _0184_ _0196_ _0232_ i_instruction[25] vssd1 vssd1 vccd1 vccd1 _0406_
+ sky130_fd_sc_hd__a32o_1
X_0821_ _0197_ _0332_ _0336_ _0337_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__a211o_1
X_0752_ _0274_ _0276_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__nand2_1
X_0683_ _0176_ i_instruction[13] _0169_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__and3b_1
X_1020_ clknet_3_0__leaf_i_clk _0049_ vssd1 vssd1 vccd1 vccd1 o_pc[2] sky130_fd_sc_hd__dfxtp_2
X_0804_ _0192_ _0215_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__nor2_1
X_0735_ _0254_ _0260_ _0209_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__a21boi_1
X_0666_ _0196_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__buf_6
X_0597_ i_stall i_flush vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__nor2_4
X_0520_ _0106_ _0099_ _0107_ vssd1 vssd1 vccd1 vccd1 o_imm_i[3] sky130_fd_sc_hd__a21oi_4
X_1003_ clknet_3_4__leaf_i_clk _0032_ vssd1 vssd1 vccd1 vccd1 o_csr_imm[1] sky130_fd_sc_hd__dfxtp_4
X_0718_ i_instruction[1] _0179_ _0224_ _0201_ _0244_ vssd1 vssd1 vccd1 vccd1 _0245_
+ sky130_fd_sc_hd__o32a_1
X_0649_ _0170_ i_instruction[8] vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__and2_4
X_0503_ _0094_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__buf_12
X_0983_ clknet_3_0__leaf_i_clk _0012_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[13] sky130_fd_sc_hd__dfxtp_2
X_0966_ _0454_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__clkbuf_1
X_0897_ _0184_ _0194_ _0404_ _0228_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__o211a_1
X_0820_ i_instruction[16] _0232_ _0228_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__a21o_1
X_0751_ i_instruction[13] _0275_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__or2_1
X_0682_ _0211_ _0183_ _0212_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__o21a_1
X_0949_ _0445_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__clkbuf_1
X_0803_ _0260_ _0302_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__or2_4
X_0734_ _0176_ i_instruction[15] i_instruction[13] _0169_ vssd1 vssd1 vccd1 vccd1
+ _0260_ sky130_fd_sc_hd__o31ai_4
X_0665_ i_instruction[0] _0180_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__nor2_8
X_0596_ _0145_ vssd1 vssd1 vccd1 vccd1 o_inst_supported sky130_fd_sc_hd__buf_2
X_1002_ clknet_3_3__leaf_i_clk _0031_ vssd1 vssd1 vccd1 vccd1 o_csr_imm[0] sky130_fd_sc_hd__dfxtp_4
X_0717_ _0179_ _0193_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__nand2_1
X_0648_ _0179_ _0180_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__nand2_4
X_0579_ o_funct3[1] o_funct3[0] _0132_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__and3b_1
X_0502_ _0092_ _0093_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__or2_1
X_0982_ clknet_3_7__leaf_i_clk _0011_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[12] sky130_fd_sc_hd__dfxtp_2
X_0965_ o_pc[13] i_pc[13] _0446_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__mux2_1
X_0896_ i_instruction[25] _0275_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__or2_1
X_0750_ _0176_ _0192_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__or2_2
X_0681_ i_instruction[15] i_instruction[13] _0169_ i_instruction[14] vssd1 vssd1 vccd1
+ vccd1 _0212_ sky130_fd_sc_hd__and4b_2
X_0948_ o_pc[5] i_pc[5] _0158_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__mux2_1
X_0879_ _0172_ i_instruction[5] _0305_ _0388_ _0181_ vssd1 vssd1 vccd1 vccd1 _0389_
+ sky130_fd_sc_hd__a311o_1
X_0802_ _0165_ o_csr_imm_sel _0319_ _0320_ _0248_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__o221a_1
X_0733_ _0187_ _0254_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__nand2_1
X_0664_ _0194_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__buf_6
X_0595_ o_inst_mret _0144_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__or2_1
X_1001_ clknet_3_3__leaf_i_clk _0030_ vssd1 vssd1 vccd1 vccd1 o_csr_imm_sel sky130_fd_sc_hd__dfxtp_4
X_0716_ _0164_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_8
X_0647_ _0171_ i_instruction[1] vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__nand2_8
X_0578_ i_flush _0079_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__nor2_8
X_0501_ instruction\[4\] _0068_ instruction\[2\] vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__and3_1
X_0981_ clknet_3_5__leaf_i_clk _0010_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[11] sky130_fd_sc_hd__dfxtp_2
X_0964_ _0453_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__clkbuf_1
X_0895_ _0398_ _0401_ _0402_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__o21a_1
X_0680_ _0169_ i_instruction[8] vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__nand2_2
X_0947_ _0444_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__clkbuf_1
X_0878_ _0177_ i_instruction[23] _0288_ i_instruction[10] _0387_ vssd1 vssd1 vccd1
+ vccd1 _0388_ sky130_fd_sc_hd__o221a_1
X_0801_ _0177_ _0233_ _0241_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__a21o_1
X_0732_ _0194_ _0255_ _0256_ _0257_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__a31o_1
X_0663_ _0193_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__buf_4
X_0594_ _0081_ o_csr_read _0141_ _0143_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__or4b_4
Xclkbuf_2_3_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_1000_ clknet_3_4__leaf_i_clk _0029_ vssd1 vssd1 vccd1 vccd1 o_funct3[1] sky130_fd_sc_hd__dfxtp_4
X_0715_ _0166_ instruction\[5\] _0167_ _0242_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__o211a_1
X_0646_ _0170_ i_instruction[0] vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__nand2_4
X_0577_ _0131_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[0] sky130_fd_sc_hd__buf_2
X_0500_ instruction\[3\] _0065_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__and2_1
X_0629_ _0163_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_0980_ clknet_3_7__leaf_i_clk _0009_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[10] sky130_fd_sc_hd__dfxtp_2
X_0963_ o_pc[12] i_pc[12] _0446_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__mux2_1
X_0894_ _0184_ _0271_ _0209_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__o21a_4
X_0946_ o_pc[4] i_pc[4] _0158_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__mux2_1
X_0877_ _0187_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__inv_2
X_0800_ _0302_ _0317_ _0318_ _0210_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__o31a_1
X_0731_ _0249_ _0221_ _0192_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__o21a_1
X_0662_ _0176_ _0192_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__nor2_2
X_0593_ _0067_ _0137_ _0142_ _0097_ valid_input vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__o311a_1
X_0929_ _0243_ o_csr_idx[9] _0309_ _0432_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__o211a_1
X_0714_ _0230_ _0231_ _0240_ _0241_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__a31o_1
X_0645_ _0172_ _0177_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__and2_4
X_0576_ o_csr_idx[5] o_csr_imm_sel _0125_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__and3_1
X_0628_ o_csr_pc_next[15] i_pc_next[15] _0158_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__mux2_1
X_0559_ o_csr_idx[7] _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 o_imm_i[27] sky130_fd_sc_hd__a21o_2
X_0962_ _0452_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__clkbuf_1
X_0893_ _0341_ _0399_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__or3_2
Xclkbuf_3_2__f_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0945_ _0443_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__clkbuf_1
X_0876_ _0210_ _0384_ _0385_ _0228_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__a211o_1
X_0730_ _0202_ _0184_ _0201_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__a21o_1
X_0661_ _0170_ _0186_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__nand2_8
X_0592_ o_csr_imm_sel o_funct3[1] o_funct3[0] _0068_ vssd1 vssd1 vccd1 vccd1 _0142_
+ sky130_fd_sc_hd__o31a_1
X_0928_ i_instruction[29] _0233_ _0402_ _0429_ _0431_ vssd1 vssd1 vccd1 vccd1 _0432_
+ sky130_fd_sc_hd__a221o_1
X_0859_ i_instruction[3] _0274_ _0196_ _0370_ _0210_ vssd1 vssd1 vccd1 vccd1 _0371_
+ sky130_fd_sc_hd__a32o_1
X_0713_ _0168_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__buf_6
X_0644_ _0176_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__buf_6
X_0575_ o_imm_i[10] _0127_ _0128_ _0130_ o_inst_branch vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[2]
+ sky130_fd_sc_hd__a311o_4
X_0627_ _0162_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__clkbuf_1
X_0558_ o_csr_idx[6] _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 o_imm_i[26] sky130_fd_sc_hd__a21o_2
X_0489_ _0085_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__buf_12
X_0961_ o_pc[11] i_pc[11] _0446_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__mux2_1
X_0892_ i_instruction[10] i_instruction[11] _0184_ _0236_ vssd1 vssd1 vccd1 vccd1
+ _0400_ sky130_fd_sc_hd__and4b_1
X_0944_ o_pc[3] i_pc[3] _0158_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__mux2_1
X_0875_ i_instruction[23] _0232_ _0196_ i_instruction[5] vssd1 vssd1 vccd1 vccd1 _0385_
+ sky130_fd_sc_hd__a22o_1
X_0660_ _0190_ _0191_ i_flush vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__a21oi_1
X_0591_ _0139_ _0140_ _0137_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__a21oi_1
X_0927_ _0228_ _0430_ i_stall vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__a21o_1
X_0858_ _0200_ _0369_ _0341_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__o21bai_1
X_0789_ _0134_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__buf_4
X_0712_ i_instruction[5] _0233_ _0239_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__a21o_1
X_0643_ i_instruction[14] vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__buf_6
X_0574_ o_csr_imm_sel o_funct3[1] _0129_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__and3b_1
X_1057_ o_csr_idx[4] vssd1 vssd1 vccd1 vccd1 o_rs2[4] sky130_fd_sc_hd__buf_2
X_0626_ o_csr_pc_next[14] i_pc_next[14] _0158_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__mux2_1
X_0557_ o_csr_idx[5] _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 o_imm_i[25] sky130_fd_sc_hd__a21o_2
X_0488_ _0064_ instruction\[3\] instruction\[2\] vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__or3b_4
X_0609_ o_csr_pc_next[6] i_pc_next[6] _0147_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__mux2_1
X_0960_ _0451_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__clkbuf_1
X_0891_ i_instruction[12] _0361_ _0260_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__a21o_1
X_0943_ _0442_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__clkbuf_1
X_0874_ _0369_ _0383_ _0341_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__o21bai_1
X_0590_ _0064_ instruction\[2\] _0074_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__a21o_1
X_0926_ _0305_ _0235_ _0194_ i_instruction[29] vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__a22o_1
X_0857_ _0221_ _0361_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__nor2_1
X_0788_ _0165_ o_funct3[0] _0307_ _0308_ _0248_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__o221a_1
X_0711_ _0186_ _0180_ _0238_ _0179_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__o22a_1
X_0642_ _0174_ instruction\[0\] vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__nand2_1
X_0573_ o_csr_idx[5] _0070_ _0128_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__o21ai_1
X_1056_ o_csr_idx[3] vssd1 vssd1 vccd1 vccd1 o_rs2[3] sky130_fd_sc_hd__buf_2
X_0909_ _0243_ o_csr_idx[6] _0309_ _0415_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__o211a_1
X_0625_ _0161_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__clkbuf_1
X_0556_ o_csr_idx[4] _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 o_imm_i[24] sky130_fd_sc_hd__a21o_2
X_0487_ _0084_ vssd1 vssd1 vccd1 vccd1 o_inst_mret sky130_fd_sc_hd__buf_2
X_1039_ o_csr_pc_next[2] vssd1 vssd1 vccd1 vccd1 o_pc_next[2] sky130_fd_sc_hd__buf_2
X_0608_ _0152_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__clkbuf_1
X_0539_ o_csr_idx[11] _0085_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__and2_1
X_0890_ _0215_ _0273_ _0333_ i_instruction[2] vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__o31a_1
X_0942_ o_pc[2] i_pc[2] _0158_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__mux2_1
X_0873_ _0172_ i_instruction[5] _0237_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__a21boi_1
X_0925_ i_instruction[10] _0215_ _0260_ _0428_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__a211o_1
X_0856_ _0166_ o_csr_idx[0] _0309_ _0368_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__o211a_1
X_0787_ i_instruction[12] _0229_ _0195_ _0168_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__a31o_1
X_0710_ _0234_ _0224_ _0237_ i_instruction[1] vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__a31oi_1
X_0641_ _0168_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__buf_4
X_0572_ instruction\[2\] _0071_ _0074_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__or3_1
X_1055_ o_csr_idx[2] vssd1 vssd1 vccd1 vccd1 o_rs2[2] sky130_fd_sc_hd__buf_2
X_0908_ _0168_ _0414_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__or2_1
X_0839_ _0295_ _0271_ _0321_ _0341_ _0180_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__o221a_1
X_0624_ o_csr_pc_next[13] i_pc_next[13] _0158_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__mux2_1
X_0555_ o_csr_idx[3] _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 o_imm_i[23] sky130_fd_sc_hd__a21o_2
X_0486_ o_csr_idx[2] o_csr_idx[1] _0083_ o_csr_idx[9] vssd1 vssd1 vccd1 vccd1 _0084_
+ sky130_fd_sc_hd__and4b_1
X_1038_ o_csr_pc_next[1] vssd1 vssd1 vccd1 vccd1 o_pc_next[1] sky130_fd_sc_hd__buf_2
Xclkbuf_3_5__f_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0607_ o_csr_pc_next[5] i_pc_next[5] _0147_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__mux2_1
X_0538_ _0092_ _0116_ _0117_ _0086_ vssd1 vssd1 vccd1 vccd1 o_imm_i[11] sky130_fd_sc_hd__o211a_2
X_0469_ instruction\[3\] instruction\[2\] _0071_ instruction\[6\] vssd1 vssd1 vccd1
+ vccd1 _0072_ sky130_fd_sc_hd__or4b_1
X_0941_ _0441_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__clkbuf_1
X_0872_ _0174_ _0381_ _0382_ _0248_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__o211a_1
X_0924_ i_instruction[12] _0178_ _0400_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__a21o_1
X_0855_ _0366_ _0367_ _0174_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__a21o_1
X_0786_ _0304_ _0306_ _0289_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__o21a_1
X_0640_ _0166_ valid_input _0167_ _0173_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__o211a_1
X_0571_ _0086_ _0127_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[4] sky130_fd_sc_hd__nand2_4
X_1054_ o_csr_idx[1] vssd1 vssd1 vccd1 vccd1 o_rs2[1] sky130_fd_sc_hd__buf_2
X_0907_ _0410_ _0412_ _0413_ _0289_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__o22a_1
X_0838_ _0174_ _0347_ _0351_ _0352_ _0134_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__o311a_1
X_0769_ _0235_ _0194_ _0291_ _0180_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__o211a_1
X_0623_ _0160_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__clkbuf_1
X_0554_ o_csr_idx[2] _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 o_imm_i[22] sky130_fd_sc_hd__a21o_2
X_0485_ _0080_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__inv_2
X_1037_ o_csr_read vssd1 vssd1 vccd1 vccd1 o_inst_csr_req sky130_fd_sc_hd__buf_2
X_0606_ _0151_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__clkbuf_1
X_0537_ o_csr_idx[0] _0068_ _0065_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__or3b_1
X_0468_ instruction\[5\] _0064_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__or2_1
X_0940_ o_pc[1] i_pc[1] _0158_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__mux2_1
X_0871_ _0164_ o_csr_idx[2] vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__or2_1
X_0923_ _0243_ o_csr_idx[8] _0309_ _0427_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__o211a_1
X_0854_ i_instruction[20] _0195_ _0273_ i_instruction[2] _0289_ vssd1 vssd1 vccd1
+ vccd1 _0367_ sky130_fd_sc_hd__a221o_1
X_0785_ i_instruction[12] _0233_ _0197_ _0305_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__a22o_1
X_0570_ o_inst_jal _0075_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__nor2_4
X_1053_ o_csr_idx[0] vssd1 vssd1 vccd1 vccd1 o_rs2[0] sky130_fd_sc_hd__buf_2
X_0906_ i_instruction[5] _0221_ _0275_ i_instruction[26] _0259_ vssd1 vssd1 vccd1
+ vccd1 _0413_ sky130_fd_sc_hd__o221a_1
X_0837_ _0164_ o_csr_imm[3] vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__or2_1
X_0768_ _0177_ _0270_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__or2_1
X_0699_ _0166_ instruction\[4\] _0167_ _0227_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__o211a_1
X_0622_ o_csr_pc_next[12] i_pc_next[12] _0158_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__mux2_1
X_0553_ o_csr_idx[1] _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 o_imm_i[21] sky130_fd_sc_hd__a21o_2
X_0484_ _0082_ vssd1 vssd1 vccd1 vccd1 o_csr_ebreak sky130_fd_sc_hd__buf_2
X_1036_ o_csr_idx[11] vssd1 vssd1 vccd1 vccd1 o_imm_i[31] sky130_fd_sc_hd__buf_2
X_0605_ o_csr_pc_next[4] i_pc_next[4] _0147_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__mux2_1
X_0536_ o_rd[0] o_csr_idx[11] _0097_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__mux2_1
X_0467_ instruction\[6\] _0069_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__or2_1
X_1019_ clknet_3_5__leaf_i_clk _0048_ vssd1 vssd1 vccd1 vccd1 o_pc[1] sky130_fd_sc_hd__dfxtp_2
X_0519_ o_rd[3] _0099_ _0086_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__o21ai_1
X_0870_ _0289_ _0377_ _0378_ _0380_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__o22a_2
X_0999_ clknet_3_3__leaf_i_clk _0028_ vssd1 vssd1 vccd1 vccd1 o_funct3[0] sky130_fd_sc_hd__dfxtp_4
X_0922_ _0425_ _0426_ _0241_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__a21o_1
X_0853_ _0197_ _0359_ _0360_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__a31o_1
X_0784_ _0187_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__buf_6
X_1052_ o_csr_pc_next[15] vssd1 vssd1 vccd1 vccd1 o_pc_next[15] sky130_fd_sc_hd__buf_2
X_0905_ i_instruction[26] _0207_ _0196_ _0411_ _0206_ vssd1 vssd1 vccd1 vccd1 _0412_
+ sky130_fd_sc_hd__a221o_1
X_0836_ i_instruction[18] _0233_ _0197_ _0348_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_
+ sky130_fd_sc_hd__a221o_1
X_0767_ i_instruction[10] _0288_ _0188_ _0250_ _0289_ vssd1 vssd1 vccd1 vccd1 _0290_
+ sky130_fd_sc_hd__a2111o_1
X_0698_ _0220_ _0226_ _0174_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__a21o_1
X_0621_ _0159_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__clkbuf_1
X_0552_ o_csr_idx[0] _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 o_imm_i[20] sky130_fd_sc_hd__a21o_2
X_0483_ o_csr_idx[0] _0081_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__and2_1
X_1035_ o_csr_imm_sel vssd1 vssd1 vccd1 vccd1 o_funct3[2] sky130_fd_sc_hd__buf_2
X_0819_ _0333_ _0335_ _0272_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__o21a_1
X_0604_ _0150_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__clkbuf_1
X_0535_ _0115_ vssd1 vssd1 vccd1 vccd1 o_imm_i[10] sky130_fd_sc_hd__clkbuf_4
X_0466_ instruction\[5\] instruction\[4\] _0063_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__nand3_1
X_1018_ clknet_3_6__leaf_i_clk _0047_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[11] sky130_fd_sc_hd__dfxtp_4
X_0518_ o_csr_idx[3] vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__inv_2
X_0998_ clknet_3_1__leaf_i_clk _0027_ vssd1 vssd1 vccd1 vccd1 o_rd[4] sky130_fd_sc_hd__dfxtp_2
X_0921_ _0305_ _0284_ _0195_ i_instruction[28] _0289_ vssd1 vssd1 vccd1 vccd1 _0426_
+ sky130_fd_sc_hd__a221o_1
X_0852_ i_instruction[20] _0232_ _0210_ _0364_ _0206_ vssd1 vssd1 vccd1 vccd1 _0365_
+ sky130_fd_sc_hd__a221o_1
X_0783_ _0299_ _0300_ _0303_ _0180_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__o31a_1
X_1051_ o_csr_pc_next[14] vssd1 vssd1 vccd1 vccd1 o_pc_next[14] sky130_fd_sc_hd__buf_2
X_0904_ i_instruction[2] _0250_ _0223_ _0249_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__a22o_1
X_0835_ _0235_ _0271_ _0349_ _0210_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__o211a_1
X_0766_ _0181_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__buf_6
X_0697_ _0221_ _0179_ _0222_ _0225_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__a31o_1
Xclkbuf_2_2_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0620_ o_csr_pc_next[11] i_pc_next[11] _0158_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__mux2_1
X_0551_ _0118_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__buf_12
X_0482_ o_csr_idx[8] _0080_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__nor2_2
X_1034_ o_alu_ctrl[3] vssd1 vssd1 vccd1 vccd1 o_csr_idx[10] sky130_fd_sc_hd__buf_2
X_0818_ i_instruction[8] _0322_ _0334_ _0321_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__a211o_1
X_0749_ _0186_ _0221_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__or2_2
X_0603_ o_csr_pc_next[3] i_pc_next[3] _0147_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__mux2_1
X_0534_ o_alu_ctrl[3] _0085_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__and2_1
X_0465_ _0068_ _0067_ vssd1 vssd1 vccd1 vccd1 o_inst_jal sky130_fd_sc_hd__nor2_4
X_1017_ clknet_3_3__leaf_i_clk _0046_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[3] sky130_fd_sc_hd__dfxtp_4
X_0517_ _0105_ vssd1 vssd1 vccd1 vccd1 o_imm_i[2] sky130_fd_sc_hd__buf_2
X_0997_ clknet_3_4__leaf_i_clk _0026_ vssd1 vssd1 vccd1 vccd1 o_rd[3] sky130_fd_sc_hd__dfxtp_2
X_0920_ i_instruction[28] _0233_ _0402_ _0424_ _0228_ vssd1 vssd1 vccd1 vccd1 _0425_
+ sky130_fd_sc_hd__a221o_1
X_0851_ _0321_ _0341_ _0362_ _0363_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__o31a_1
X_0782_ i_instruction[13] _0273_ _0236_ _0301_ _0302_ vssd1 vssd1 vccd1 vccd1 _0303_
+ sky130_fd_sc_hd__a221o_1
X_1050_ o_csr_pc_next[13] vssd1 vssd1 vccd1 vccd1 o_pc_next[13] sky130_fd_sc_hd__buf_2
X_0903_ _0401_ _0408_ _0409_ _0402_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__o31a_1
X_0834_ _0291_ _0274_ _0302_ _0341_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__a211o_1
X_0765_ _0171_ _0186_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__and2_1
X_0696_ i_instruction[4] _0207_ _0210_ _0224_ _0206_ vssd1 vssd1 vccd1 vccd1 _0225_
+ sky130_fd_sc_hd__a221o_1
X_0550_ _0093_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__buf_12
X_0481_ o_csr_imm_sel o_funct3[1] o_funct3[0] _0079_ vssd1 vssd1 vccd1 vccd1 _0080_
+ sky130_fd_sc_hd__or4_1
X_1033_ clknet_3_2__leaf_i_clk _0062_ vssd1 vssd1 vccd1 vccd1 o_pc[15] sky130_fd_sc_hd__dfxtp_2
X_0817_ _0171_ i_instruction[6] _0212_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__and3_1
X_0748_ _0223_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__buf_4
X_0679_ _0209_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__buf_4
X_0602_ _0149_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__clkbuf_1
X_0533_ _0114_ vssd1 vssd1 vccd1 vccd1 o_imm_i[9] sky130_fd_sc_hd__buf_2
X_0464_ instruction\[3\] vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkinv_2
X_1016_ clknet_3_6__leaf_i_clk _0045_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[9] sky130_fd_sc_hd__dfxtp_4
X_0516_ _0086_ _0104_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__and2_1
X_0996_ clknet_3_6__leaf_i_clk _0025_ vssd1 vssd1 vccd1 vccd1 o_rd[2] sky130_fd_sc_hd__dfxtp_2
X_0850_ _0199_ _0260_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__nand2_1
X_0781_ _0176_ i_instruction[13] _0169_ i_instruction[12] vssd1 vssd1 vccd1 vccd1
+ _0302_ sky130_fd_sc_hd__and4b_2
X_0979_ clknet_3_7__leaf_i_clk _0008_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[9] sky130_fd_sc_hd__dfxtp_2
X_0902_ _0249_ _0215_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__and2_1
X_0833_ _0305_ _0235_ _0325_ i_instruction[10] vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__a22o_1
X_0764_ _0165_ o_rd[2] _0282_ _0287_ _0248_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__o221a_1
X_0695_ _0215_ _0223_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__nor2_4
X_0480_ instruction\[6\] _0078_ _0076_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__nand3_4
X_1032_ clknet_3_5__leaf_i_clk _0061_ vssd1 vssd1 vccd1 vccd1 o_pc[14] sky130_fd_sc_hd__dfxtp_2
X_0816_ _0211_ _0183_ _0212_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__nor3b_4
X_0747_ _0182_ _0271_ _0209_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__o21a_1
X_0678_ i_instruction[1] _0179_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__nor2_4
X_0601_ o_csr_pc_next[2] i_pc_next[2] _0147_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__mux2_1
X_0532_ o_csr_idx[9] _0085_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__and2_1
X_0463_ instruction\[3\] _0067_ vssd1 vssd1 vccd1 vccd1 o_inst_jalr sky130_fd_sc_hd__nor2_4
X_1015_ clknet_3_6__leaf_i_clk _0044_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[8] sky130_fd_sc_hd__dfxtp_4
X_0515_ o_rd[2] o_csr_idx[2] _0099_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__mux2_1
X_0995_ clknet_3_4__leaf_i_clk _0024_ vssd1 vssd1 vccd1 vccd1 o_rd[1] sky130_fd_sc_hd__dfxtp_2
X_0780_ i_instruction[11] _0235_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__nand2_2
X_0978_ clknet_3_0__leaf_i_clk _0007_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[8] sky130_fd_sc_hd__dfxtp_2
X_0901_ _0223_ _0333_ i_instruction[5] vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__o21a_1
X_0832_ i_instruction[18] _0178_ _0315_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__o21a_1
X_0763_ i_instruction[9] _0283_ _0285_ _0286_ _0168_ vssd1 vssd1 vccd1 vccd1 _0287_
+ sky130_fd_sc_hd__a221o_1
X_0694_ _0170_ _0176_ _0186_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__and3_4
X_1031_ clknet_3_2__leaf_i_clk _0060_ vssd1 vssd1 vccd1 vccd1 o_pc[13] sky130_fd_sc_hd__dfxtp_2
X_0815_ _0182_ _0331_ _0178_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__a21o_1
X_0746_ _0187_ _0270_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__nand2_2
X_0677_ _0206_ _0193_ _0207_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__a21o_4
X_0600_ _0148_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__clkbuf_1
X_0531_ _0113_ vssd1 vssd1 vccd1 vccd1 o_imm_i[8] sky130_fd_sc_hd__buf_2
Xclkbuf_3_1__f_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0462_ instruction\[2\] _0065_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__nand2_4
X_1014_ clknet_3_4__leaf_i_clk _0043_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[7] sky130_fd_sc_hd__dfxtp_2
X_0729_ _0254_ _0201_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__nand2_1
X_0514_ _0103_ vssd1 vssd1 vccd1 vccd1 o_imm_i[1] sky130_fd_sc_hd__buf_2
X_0994_ clknet_3_1__leaf_i_clk _0023_ vssd1 vssd1 vccd1 vccd1 o_rd[0] sky130_fd_sc_hd__dfxtp_4
X_0977_ clknet_3_2__leaf_i_clk _0006_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[7] sky130_fd_sc_hd__dfxtp_2
X_0900_ _0243_ o_csr_idx[5] _0309_ _0407_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__o211a_1
X_0831_ _0165_ o_csr_imm[2] _0344_ _0346_ _0248_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__o221a_1
X_0762_ i_instruction[4] _0273_ _0277_ i_instruction[9] _0260_ vssd1 vssd1 vccd1 vccd1
+ _0286_ sky130_fd_sc_hd__a221o_1
X_0693_ _0192_ _0201_ _0204_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__or3_1
X_1030_ clknet_3_5__leaf_i_clk _0059_ vssd1 vssd1 vccd1 vccd1 o_pc[12] sky130_fd_sc_hd__dfxtp_2
X_0814_ _0192_ _0184_ _0201_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__or3b_4
X_0745_ _0171_ i_instruction[13] vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__nand2_1
X_0676_ _0179_ _0180_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__nor2_2
X_0530_ o_csr_idx[8] _0085_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__and2_1
X_0461_ _0066_ vssd1 vssd1 vccd1 vccd1 o_inst_branch sky130_fd_sc_hd__clkbuf_4
X_1013_ clknet_3_6__leaf_i_clk _0042_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[6] sky130_fd_sc_hd__dfxtp_4
X_0728_ _0171_ _0249_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__nand2_1
X_0659_ _0174_ instruction\[1\] vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__nand2_1
X_0513_ _0086_ _0102_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__and2_1
X_0993_ clknet_3_1__leaf_i_clk _0022_ vssd1 vssd1 vccd1 vccd1 instruction\[6\] sky130_fd_sc_hd__dfxtp_4
X_0976_ clknet_3_0__leaf_i_clk _0005_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[6] sky130_fd_sc_hd__dfxtp_2
X_0830_ _0229_ _0345_ _0241_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__a21o_1
X_0761_ _0284_ _0271_ _0209_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__o21a_1
X_0692_ _0170_ _0176_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__nand2_8
X_0959_ o_pc[10] i_pc[10] _0446_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__mux2_1
X_0813_ _0177_ _0182_ _0195_ i_instruction[16] _0189_ vssd1 vssd1 vccd1 vccd1 _0330_
+ sky130_fd_sc_hd__a221o_1
X_0744_ i_instruction[8] _0194_ _0250_ i_instruction[3] _0268_ vssd1 vssd1 vccd1 vccd1
+ _0269_ sky130_fd_sc_hd__a221o_1
X_0675_ _0179_ _0180_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__and2_2
X_0460_ _0063_ _0065_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__and2_1
X_1012_ clknet_3_4__leaf_i_clk _0041_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[5] sky130_fd_sc_hd__dfxtp_4
X_0727_ _0249_ _0194_ _0250_ i_instruction[2] _0252_ vssd1 vssd1 vccd1 vccd1 _0253_
+ sky130_fd_sc_hd__a221o_1
X_0658_ _0175_ _0190_ i_flush vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a21oi_1
X_0589_ instruction\[6\] _0138_ instruction\[4\] instruction\[2\] vssd1 vssd1 vccd1
+ vccd1 _0139_ sky130_fd_sc_hd__or4b_1
X_0512_ o_rd[1] o_csr_idx[1] _0099_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__mux2_4
X_0992_ clknet_3_1__leaf_i_clk _0021_ vssd1 vssd1 vccd1 vccd1 instruction\[5\] sky130_fd_sc_hd__dfxtp_4
X_0975_ clknet_3_7__leaf_i_clk _0004_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[5] sky130_fd_sc_hd__dfxtp_2
X_0760_ _0172_ i_instruction[9] vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__and2_2
X_0691_ i_instruction[4] _0195_ _0189_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__a21o_1
X_0958_ _0450_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__clkbuf_1
X_0889_ _0243_ o_csr_idx[4] _0309_ _0397_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__o211a_1
X_0812_ _0165_ o_csr_imm[0] _0324_ _0329_ _0248_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__o221a_1
X_0743_ _0251_ _0200_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__nor2_1
X_0674_ _0201_ _0204_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__nor2_1
X_1011_ clknet_3_4__leaf_i_clk _0040_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[4] sky130_fd_sc_hd__dfxtp_4
X_0726_ _0251_ _0199_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__nor2_1
X_0657_ _0178_ _0189_ _0165_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__o21ai_2
X_0588_ o_csr_imm_sel o_funct3[1] instruction\[5\] _0068_ vssd1 vssd1 vccd1 vccd1
+ _0138_ sky130_fd_sc_hd__or4_1
X_0511_ _0101_ vssd1 vssd1 vccd1 vccd1 o_imm_i[0] sky130_fd_sc_hd__buf_2
X_0709_ i_instruction[11] _0235_ _0236_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__nand3_2
X_0991_ clknet_3_1__leaf_i_clk _0020_ vssd1 vssd1 vccd1 vccd1 instruction\[4\] sky130_fd_sc_hd__dfxtp_2
X_0974_ clknet_3_2__leaf_i_clk _0003_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[4] sky130_fd_sc_hd__dfxtp_2
X_0690_ _0166_ instruction\[3\] _0167_ _0219_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__o211a_1
Xclkbuf_3_4__f_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0957_ o_pc[9] i_pc[9] _0446_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__mux2_1
X_0888_ _0210_ _0393_ _0396_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__a21o_1
X_0811_ _0197_ _0259_ _0326_ _0328_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__a31o_1
X_0742_ i_instruction[1] _0182_ _0266_ _0168_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__a31o_1
X_0673_ _0202_ _0203_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__nor2_1
X_1010_ clknet_3_4__leaf_i_clk _0039_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[3] sky130_fd_sc_hd__dfxtp_4
X_0725_ _0188_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__inv_2
X_0656_ _0181_ _0188_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__or2_1
X_0587_ instruction\[5\] _0064_ _0063_ _0137_ vssd1 vssd1 vccd1 vccd1 o_reg_write
+ sky130_fd_sc_hd__a31oi_4
X_0510_ _0095_ _0100_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__and2b_2
X_0708_ i_instruction[14] i_instruction[13] i_instruction[15] i_ready vssd1 vssd1
+ vccd1 vccd1 _0236_ sky130_fd_sc_hd__and4bb_4
X_0639_ _0168_ _0172_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__or2_1
X_0990_ clknet_3_1__leaf_i_clk _0019_ vssd1 vssd1 vccd1 vccd1 instruction\[3\] sky130_fd_sc_hd__dfxtp_4
X_0973_ clknet_3_0__leaf_i_clk _0002_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[3] sky130_fd_sc_hd__dfxtp_2
X_0956_ _0449_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__clkbuf_1
X_0887_ _0172_ _0229_ _0394_ _0395_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__a31o_1
X_0810_ _0186_ _0233_ _0327_ i_stall vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__a211o_1
X_0741_ _0221_ _0201_ _0192_ i_instruction[0] vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__a211o_1
X_0672_ _0171_ i_instruction[12] vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__nand2_2
X_0939_ o_csr_idx[11] _0243_ _0439_ _0440_ _0167_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__o221a_1
X_0724_ _0186_ _0221_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__nor2_2
X_0655_ _0182_ _0183_ _0184_ _0185_ _0187_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__o41a_2
X_0586_ instruction\[1\] instruction\[0\] vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__nand2_2
X_0707_ _0171_ i_instruction[10] vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__and2_4
X_0638_ _0171_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__buf_4
X_0569_ _0126_ vssd1 vssd1 vccd1 vccd1 o_alu_ctrl[1] sky130_fd_sc_hd__buf_2
X_0972_ clknet_3_6__leaf_i_clk _0001_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[2] sky130_fd_sc_hd__dfxtp_2
X_0955_ o_pc[8] i_pc[8] _0446_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__mux2_1
X_0886_ i_instruction[24] _0232_ _0196_ i_instruction[6] i_stall vssd1 vssd1 vccd1
+ vccd1 _0395_ sky130_fd_sc_hd__a221o_1
X_0740_ _0166_ o_rd[0] _0167_ _0265_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__o211a_1
X_0671_ _0182_ _0183_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__or2_2
X_0938_ i_instruction[31] _0208_ _0241_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__a21o_1
X_0869_ _0341_ _0379_ _0210_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__o21a_1
Xclkbuf_2_1_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0723_ i_instruction[7] vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__buf_4
X_0654_ _0176_ _0186_ _0170_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__o21ai_4
X_0585_ _0136_ vssd1 vssd1 vccd1 vccd1 o_csr_clear sky130_fd_sc_hd__buf_2
X_0706_ _0211_ _0183_ _0212_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__o21ai_4
X_0637_ _0170_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__buf_6
X_0568_ o_csr_idx[5] _0125_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__and2_1
X_0499_ _0091_ vssd1 vssd1 vccd1 vccd1 o_rs1[4] sky130_fd_sc_hd__buf_2
X_0971_ clknet_3_2__leaf_i_clk _0000_ vssd1 vssd1 vccd1 vccd1 o_csr_pc_next[1] sky130_fd_sc_hd__dfxtp_2
X_0954_ _0448_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__clkbuf_1
X_0885_ i_instruction[11] _0192_ _0194_ i_instruction[24] vssd1 vssd1 vccd1 vccd1
+ _0394_ sky130_fd_sc_hd__a22o_1
X_0670_ _0185_ _0198_ _0199_ _0200_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__nand4b_4
X_0937_ _0321_ _0428_ _0402_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__o21a_1
X_0868_ _0198_ _0369_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__nor2_1
X_0799_ _0185_ _0301_ _0236_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__o21a_1
X_0722_ _0243_ instruction\[6\] _0246_ _0247_ _0248_ vssd1 vssd1 vccd1 vccd1 _0022_
+ sky130_fd_sc_hd__o221a_1
X_0653_ i_instruction[15] vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__buf_6
X_0584_ o_funct3[1] o_funct3[0] _0132_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__and3_1
X_0705_ _0232_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__buf_6
X_0636_ _0169_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__buf_8
X_0567_ instruction\[6\] _0069_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__nor2_1
X_0498_ o_csr_imm[4] _0085_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__and2_1
Xclkbuf_3_7__f_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0619_ _0146_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__buf_12
X_0970_ _0456_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__clkbuf_1
X_0953_ o_pc[7] i_pc[7] _0446_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__mux2_1
X_0884_ _0172_ i_instruction[6] _0391_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__a31o_1
X_0936_ _0165_ o_alu_ctrl[3] _0437_ _0438_ _0167_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__o221a_1
X_0867_ i_instruction[22] _0232_ _0197_ i_instruction[4] _0228_ vssd1 vssd1 vccd1
+ vccd1 _0378_ sky130_fd_sc_hd__a221o_1
X_0798_ _0234_ _0198_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__nor2_1
X_0721_ _0134_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__buf_6
X_0652_ i_instruction[5] i_instruction[6] _0169_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__o21a_1
X_0583_ _0135_ vssd1 vssd1 vccd1 vccd1 o_csr_set sky130_fd_sc_hd__buf_2
X_0919_ i_instruction[4] _0333_ _0401_ _0423_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__a211o_1
X_0704_ _0207_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_8
X_0635_ i_ready vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__buf_4
X_0566_ _0092_ _0124_ instruction\[2\] vssd1 vssd1 vccd1 vccd1 o_op1_src sky130_fd_sc_hd__o21a_2
X_0497_ _0090_ vssd1 vssd1 vccd1 vccd1 o_rs1[3] sky130_fd_sc_hd__buf_2
X_1049_ o_csr_pc_next[12] vssd1 vssd1 vccd1 vccd1 o_pc_next[12] sky130_fd_sc_hd__buf_2
X_0618_ _0157_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__clkbuf_1
X_0549_ o_csr_imm[4] _0095_ _0120_ vssd1 vssd1 vccd1 vccd1 o_imm_i[19] sky130_fd_sc_hd__a21o_2
X_0952_ _0447_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__clkbuf_1
X_0883_ i_instruction[11] _0215_ _0333_ i_instruction[6] _0341_ vssd1 vssd1 vccd1
+ vccd1 _0392_ sky130_fd_sc_hd__a221o_1
X_0935_ i_instruction[30] _0208_ _0241_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__a21o_1
X_0866_ i_instruction[22] _0194_ _0273_ i_instruction[4] _0376_ vssd1 vssd1 vccd1
+ vccd1 _0377_ sky130_fd_sc_hd__a221o_1
X_0797_ _0166_ o_funct3[1] _0309_ _0316_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__o211a_1
X_0720_ i_instruction[6] _0208_ _0241_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__a21o_1
X_0651_ _0169_ i_instruction[12] vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__and2_4
X_0582_ o_funct3[0] _0134_ _0123_ o_funct3[1] vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__and4b_1
X_0918_ i_instruction[9] _0215_ _0223_ i_instruction[12] vssd1 vssd1 vccd1 vccd1 _0423_
+ sky130_fd_sc_hd__a22o_1
X_0849_ _0236_ _0361_ _0199_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__o21ba_1
X_0703_ i_instruction[5] _0177_ _0181_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__or3_1
X_0634_ i_stall vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__buf_6
X_0565_ _0071_ _0074_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__nor2_1
X_0496_ o_csr_imm[3] _0086_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__and2_1
X_1048_ o_csr_pc_next[11] vssd1 vssd1 vccd1 vccd1 o_pc_next[11] sky130_fd_sc_hd__buf_2
X_0617_ o_csr_pc_next[10] i_pc_next[10] _0147_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__mux2_1
X_0548_ o_csr_imm[3] _0095_ _0120_ vssd1 vssd1 vccd1 vccd1 o_imm_i[18] sky130_fd_sc_hd__a21o_2
X_0479_ instruction\[5\] instruction\[4\] _0063_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__and3_1
X_0951_ o_pc[6] i_pc[6] _0446_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__mux2_1
X_0882_ _0236_ _0301_ _0260_ _0361_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__a211o_1
X_0934_ _0435_ _0436_ _0402_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__o21a_1
X_0865_ _0186_ _0375_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__nor2_1
X_0796_ _0289_ _0314_ _0315_ _0276_ _0168_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__a221o_1
X_0650_ i_instruction[7] i_instruction[9] i_instruction[10] i_instruction[11] _0169_
+ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__o41a_4
X_0581_ i_flush vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__clkinv_2
X_0917_ _0174_ _0421_ _0422_ _0248_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__o211a_1
X_0848_ i_instruction[15] i_instruction[13] _0169_ _0176_ vssd1 vssd1 vccd1 vccd1
+ _0361_ sky130_fd_sc_hd__and4bb_2
X_0779_ _0172_ i_instruction[5] i_instruction[6] _0236_ vssd1 vssd1 vccd1 vccd1 _0300_
+ sky130_fd_sc_hd__and4_1
X_0702_ _0229_ _0192_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__nand2_1
X_0633_ _0134_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_8
X_0564_ o_csr_imm_sel o_funct3[1] o_funct3[0] _0123_ vssd1 vssd1 vccd1 vccd1 o_csr_read
+ sky130_fd_sc_hd__o31a_4
X_0495_ _0089_ vssd1 vssd1 vccd1 vccd1 o_rs1[2] sky130_fd_sc_hd__buf_2
X_1047_ o_csr_pc_next[10] vssd1 vssd1 vccd1 vccd1 o_pc_next[10] sky130_fd_sc_hd__buf_2
X_0616_ _0156_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__clkbuf_1
X_0547_ o_csr_imm[2] _0095_ _0120_ vssd1 vssd1 vccd1 vccd1 o_imm_i[17] sky130_fd_sc_hd__a21o_2
X_0478_ o_res_src[1] o_res_src[2] vssd1 vssd1 vccd1 vccd1 o_res_src[0] sky130_fd_sc_hd__nor2_4
X_0950_ _0146_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__buf_12
X_0881_ _0243_ o_csr_idx[3] _0309_ _0390_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__o211a_1
Xclkbuf_3_0__f_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0933_ i_instruction[12] _0178_ _0215_ i_instruction[8] _0260_ vssd1 vssd1 vccd1
+ vccd1 _0436_ sky130_fd_sc_hd__a221o_1
X_0864_ _0172_ i_instruction[6] vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__nand2_1
X_0795_ _0181_ _0187_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__nor2_2
X_0580_ _0133_ vssd1 vssd1 vccd1 vccd1 o_csr_write sky130_fd_sc_hd__buf_2
X_0916_ _0164_ o_csr_idx[7] vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__or2_1
X_0847_ _0305_ _0199_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__nand2_1
X_0778_ _0234_ _0199_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__nor2_1
X_0701_ _0228_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__buf_6
X_0632_ _0165_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_8
X_0563_ instruction\[6\] _0078_ _0076_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__and3_1
X_0494_ o_csr_imm[2] _0086_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__and2_1
X_1046_ o_csr_pc_next[9] vssd1 vssd1 vccd1 vccd1 o_pc_next[9] sky130_fd_sc_hd__buf_2
X_0615_ o_csr_pc_next[9] i_pc_next[9] _0147_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__mux2_1
X_0546_ o_csr_imm[1] _0095_ _0120_ vssd1 vssd1 vccd1 vccd1 o_imm_i[16] sky130_fd_sc_hd__a21o_2
X_0477_ _0067_ vssd1 vssd1 vccd1 vccd1 o_res_src[1] sky130_fd_sc_hd__clkinv_4
X_1029_ clknet_3_0__leaf_i_clk _0058_ vssd1 vssd1 vccd1 vccd1 o_pc[11] sky130_fd_sc_hd__dfxtp_2
X_0529_ _0112_ vssd1 vssd1 vccd1 vccd1 o_imm_i[7] sky130_fd_sc_hd__buf_2
X_0880_ _0386_ _0389_ _0241_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__a21o_1
X_0932_ _0235_ _0295_ _0236_ _0434_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__o211a_1
X_0863_ _0243_ o_csr_idx[1] _0309_ _0374_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__o211a_1
X_0794_ i_instruction[13] _0232_ _0196_ _0177_ _0313_ vssd1 vssd1 vccd1 vccd1 _0314_
+ sky130_fd_sc_hd__a221o_1
X_0915_ _0417_ _0419_ _0420_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__o21a_1
X_0846_ i_instruction[2] _0273_ _0358_ _0193_ _0305_ vssd1 vssd1 vccd1 vccd1 _0359_
+ sky130_fd_sc_hd__a221o_1
X_0777_ _0174_ _0297_ _0298_ _0248_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__o211a_1
X_0700_ _0206_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__buf_4
X_0631_ _0164_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__buf_6
X_0562_ o_alu_ctrl[3] _0093_ _0118_ vssd1 vssd1 vccd1 vccd1 o_imm_i[30] sky130_fd_sc_hd__a21o_2
X_0493_ _0088_ vssd1 vssd1 vccd1 vccd1 o_rs1[1] sky130_fd_sc_hd__buf_2
X_1045_ o_csr_pc_next[8] vssd1 vssd1 vccd1 vccd1 o_pc_next[8] sky130_fd_sc_hd__buf_2
X_0829_ _0177_ _0284_ _0195_ i_instruction[17] vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__a22o_1
X_0614_ _0155_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__clkbuf_1
X_0545_ o_csr_imm[0] _0095_ _0120_ vssd1 vssd1 vccd1 vccd1 o_imm_i[15] sky130_fd_sc_hd__a21o_2
X_0476_ _0077_ vssd1 vssd1 vccd1 vccd1 o_res_src[2] sky130_fd_sc_hd__clkbuf_4
X_1028_ clknet_3_5__leaf_i_clk _0057_ vssd1 vssd1 vccd1 vccd1 o_pc[10] sky130_fd_sc_hd__dfxtp_2
X_0528_ o_csr_idx[7] _0085_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__and2_2
X_0459_ instruction\[6\] instruction\[5\] _0064_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__and3_1
X_0931_ _0185_ _0301_ _0433_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__o21ai_1
X_0862_ _0372_ _0373_ _0241_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__a21o_1
X_0793_ _0302_ _0310_ _0312_ _0180_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__o31a_1
X_0914_ _0305_ _0182_ _0195_ i_instruction[27] _0181_ vssd1 vssd1 vccd1 vccd1 _0420_
+ sky130_fd_sc_hd__a221o_1
X_0845_ _0202_ _0203_ _0201_ _0199_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__o31ai_1
X_0776_ _0165_ o_rd[4] vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__or2_1
X_0630_ i_stall vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__inv_2
X_0561_ o_csr_idx[9] _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 o_imm_i[29] sky130_fd_sc_hd__a21o_2
X_0492_ o_csr_imm[1] _0086_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__and2_1
X_1044_ o_csr_pc_next[7] vssd1 vssd1 vccd1 vccd1 o_pc_next[7] sky130_fd_sc_hd__buf_2
X_0828_ i_instruction[17] _0233_ _0197_ _0340_ _0343_ vssd1 vssd1 vccd1 vccd1 _0344_
+ sky130_fd_sc_hd__a221o_1
X_0759_ _0244_ _0201_ _0180_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__o21ba_2
X_0613_ o_csr_pc_next[8] i_pc_next[8] _0147_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__mux2_1
X_0544_ o_csr_imm_sel _0095_ _0120_ vssd1 vssd1 vccd1 vccd1 o_imm_i[14] sky130_fd_sc_hd__a21o_2
X_0475_ instruction\[5\] _0075_ _0076_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__and3b_1
X_1027_ clknet_3_7__leaf_i_clk _0056_ vssd1 vssd1 vccd1 vccd1 o_pc[9] sky130_fd_sc_hd__dfxtp_2
X_0527_ _0111_ vssd1 vssd1 vccd1 vccd1 o_imm_i[6] sky130_fd_sc_hd__buf_2
X_0458_ instruction\[4\] vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__clkinv_2
X_0930_ i_instruction[10] _0203_ _0295_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__o21a_1
X_0861_ i_instruction[21] _0195_ _0273_ i_instruction[3] _0289_ vssd1 vssd1 vccd1
+ vccd1 _0373_ sky130_fd_sc_hd__a221o_1
X_0792_ i_instruction[6] _0311_ _0236_ i_instruction[11] vssd1 vssd1 vccd1 vccd1 _0312_
+ sky130_fd_sc_hd__o211a_1
X_0913_ i_instruction[27] _0232_ _0197_ _0418_ _0228_ vssd1 vssd1 vccd1 vccd1 _0419_
+ sky130_fd_sc_hd__a221o_1
X_0844_ _0165_ o_csr_imm[4] _0356_ _0357_ _0167_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__o221a_1
X_0775_ _0186_ _0289_ _0295_ _0296_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__o211a_1
X_0560_ o_csr_idx[8] _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 o_imm_i[28] sky130_fd_sc_hd__a21o_2
X_0491_ _0087_ vssd1 vssd1 vccd1 vccd1 o_rs1[0] sky130_fd_sc_hd__buf_2
X_1043_ o_csr_pc_next[6] vssd1 vssd1 vccd1 vccd1 o_pc_next[6] sky130_fd_sc_hd__buf_2
X_0827_ _0321_ _0341_ _0342_ _0285_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__o31a_1
X_0758_ _0280_ _0281_ _0229_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__o21a_1
X_0689_ i_instruction[3] _0208_ _0216_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a21o_1
X_0612_ _0154_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__clkbuf_1
X_0543_ o_funct3[1] _0095_ _0120_ vssd1 vssd1 vccd1 vccd1 o_imm_i[13] sky130_fd_sc_hd__a21o_2
X_0474_ instruction\[1\] instruction\[0\] vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__and2_2
X_1026_ clknet_3_0__leaf_i_clk _0055_ vssd1 vssd1 vccd1 vccd1 o_pc[8] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_3_3__f_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0526_ o_csr_idx[6] _0085_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__and2_1
X_0457_ instruction\[3\] instruction\[2\] vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__nor2_2
X_1009_ clknet_3_4__leaf_i_clk _0038_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[2] sky130_fd_sc_hd__dfxtp_4
X_0509_ o_rd[0] o_inst_store _0099_ o_csr_idx[0] vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__a22o_1
X_0860_ i_instruction[21] _0233_ _0371_ _0229_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__a211o_1
X_0791_ _0171_ i_instruction[10] vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__nand2_1
X_0989_ clknet_3_1__leaf_i_clk _0018_ vssd1 vssd1 vccd1 vccd1 instruction\[2\] sky130_fd_sc_hd__dfxtp_4
X_0912_ i_instruction[3] _0250_ _0273_ i_instruction[8] vssd1 vssd1 vccd1 vccd1 _0418_
+ sky130_fd_sc_hd__a22o_1
X_0843_ i_instruction[19] _0229_ _0195_ _0168_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__a31o_1
X_0774_ _0177_ _0228_ _0260_ _0283_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__or4_1
Xclkbuf_2_0_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_0490_ o_csr_imm[0] _0086_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__and2_1
X_1042_ o_csr_pc_next[5] vssd1 vssd1 vccd1 vccd1 o_pc_next[5] sky130_fd_sc_hd__buf_2
X_0826_ i_instruction[9] _0322_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__and2_1
X_0757_ i_instruction[9] _0194_ _0273_ i_instruction[6] vssd1 vssd1 vccd1 vccd1 _0281_
+ sky130_fd_sc_hd__a22o_1
X_0688_ _0166_ instruction\[2\] _0167_ _0218_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__o211a_1
X_0611_ o_csr_pc_next[7] i_pc_next[7] _0147_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__mux2_1
X_0542_ o_funct3[0] _0095_ _0120_ vssd1 vssd1 vccd1 vccd1 o_imm_i[12] sky130_fd_sc_hd__a21o_2
X_0473_ instruction\[4\] _0074_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__nor2_2
X_1025_ clknet_3_5__leaf_i_clk _0054_ vssd1 vssd1 vccd1 vccd1 o_pc[7] sky130_fd_sc_hd__dfxtp_2
X_0809_ _0249_ _0221_ _0315_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__o21a_1
X_0525_ _0110_ vssd1 vssd1 vccd1 vccd1 o_imm_i[5] sky130_fd_sc_hd__buf_2
X_1008_ clknet_3_4__leaf_i_clk _0037_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[1] sky130_fd_sc_hd__dfxtp_4
X_0508_ _0098_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__buf_8
X_0790_ _0234_ _0200_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__nor2_1
X_0988_ clknet_3_1__leaf_i_clk _0017_ vssd1 vssd1 vccd1 vccd1 instruction\[1\] sky130_fd_sc_hd__dfxtp_1
X_0911_ _0401_ _0416_ _0402_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__o21a_1
X_0842_ _0353_ _0355_ _0289_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__o21a_1
X_0773_ _0171_ i_instruction[11] vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__and2_1
X_1041_ o_csr_pc_next[4] vssd1 vssd1 vccd1 vccd1 o_pc_next[4] sky130_fd_sc_hd__buf_2
X_0825_ _0211_ _0183_ _0184_ _0212_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__o211a_4
X_0756_ _0251_ _0274_ _0198_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__a21oi_1
X_0687_ _0195_ _0197_ _0205_ _0217_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__a31o_1
X_0610_ _0153_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__clkbuf_1
X_0541_ _0119_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__buf_12
X_0472_ instruction\[6\] instruction\[3\] vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__or2_2
X_1024_ clknet_3_0__leaf_i_clk _0053_ vssd1 vssd1 vccd1 vccd1 o_pc[6] sky130_fd_sc_hd__dfxtp_2
X_0808_ _0249_ _0325_ _0305_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__a21o_1
X_0739_ _0229_ _0253_ _0264_ _0241_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__a211o_1
X_0524_ o_csr_idx[5] _0085_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__and2_1
X_1007_ clknet_3_4__leaf_i_clk _0036_ vssd1 vssd1 vccd1 vccd1 o_csr_idx[0] sky130_fd_sc_hd__dfxtp_4
X_0507_ _0096_ _0097_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__and2_1
X_0987_ clknet_3_1__leaf_i_clk _0016_ vssd1 vssd1 vccd1 vccd1 instruction\[0\] sky130_fd_sc_hd__dfxtp_1
X_0910_ _0375_ _0224_ _0333_ i_instruction[3] vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__a2bb2o_1
X_0841_ i_instruction[19] _0233_ _0331_ _0354_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__a22o_1
X_0772_ _0166_ o_rd[3] _0167_ _0294_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__o211a_1
X_1040_ o_csr_pc_next[3] vssd1 vssd1 vccd1 vccd1 o_pc_next[3] sky130_fd_sc_hd__buf_2
X_0824_ _0305_ _0284_ _0325_ i_instruction[9] vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__a22o_1
X_0755_ _0243_ o_rd[1] _0267_ _0279_ _0248_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__o221a_1
X_0686_ i_instruction[2] _0208_ _0210_ _0213_ _0216_ vssd1 vssd1 vccd1 vccd1 _0217_
+ sky130_fd_sc_hd__a221o_1
X_0540_ _0092_ _0118_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__and2b_1
X_0471_ _0073_ vssd1 vssd1 vccd1 vccd1 o_op2_src sky130_fd_sc_hd__buf_2
X_1023_ clknet_3_5__leaf_i_clk _0052_ vssd1 vssd1 vccd1 vccd1 o_pc[5] sky130_fd_sc_hd__dfxtp_2
X_0807_ _0203_ _0201_ _0275_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__a21oi_2
X_0738_ _0197_ _0258_ _0259_ _0263_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__a31o_1
X_0669_ _0170_ i_instruction[3] vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__nand2_4
X_0523_ _0108_ _0099_ _0109_ vssd1 vssd1 vccd1 vccd1 o_imm_i[4] sky130_fd_sc_hd__a21oi_4
X_1006_ clknet_3_6__leaf_i_clk _0035_ vssd1 vssd1 vccd1 vccd1 o_csr_imm[4] sky130_fd_sc_hd__dfxtp_4
X_0506_ o_inst_branch _0076_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__nand2_1
X_0986_ clknet_3_1__leaf_i_clk _0015_ vssd1 vssd1 vccd1 vccd1 valid_input sky130_fd_sc_hd__dfxtp_1
X_0840_ i_instruction[11] _0221_ _0196_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__and3_1
X_0771_ _0290_ _0293_ _0174_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__a21o_1
X_0969_ o_pc[15] i_pc[15] _0446_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6__f_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_0823_ _0166_ o_csr_imm[1] _0309_ _0339_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__o211a_1
X_0754_ _0229_ _0269_ _0272_ _0278_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__a22o_1
X_0685_ _0210_ _0215_ i_stall vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__a21o_1
X_0470_ o_inst_branch _0070_ _0072_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__and3b_1
X_1022_ clknet_3_2__leaf_i_clk _0051_ vssd1 vssd1 vccd1 vccd1 o_pc[4] sky130_fd_sc_hd__dfxtp_2
X_0806_ _0321_ _0323_ _0261_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__o21a_1
X_0737_ _0249_ _0232_ _0261_ _0262_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__a22o_1
X_0668_ _0170_ i_instruction[2] vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__nand2_4
X_0599_ o_csr_pc_next[1] i_pc_next[1] _0147_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__mux2_1
X_0522_ o_rd[4] _0099_ _0086_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__o21ai_1
X_1005_ clknet_3_1__leaf_i_clk _0034_ vssd1 vssd1 vccd1 vccd1 o_csr_imm[3] sky130_fd_sc_hd__dfxtp_2
X_0505_ _0096_ vssd1 vssd1 vccd1 vccd1 o_inst_store sky130_fd_sc_hd__inv_2
.ends

