** sch_path: /media/FlexRV32/asic/blocks/rom/rom_dec.sch
**.subckt rom_dec A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2]
*+ ROW[255],ROW[254],ROW[253],ROW[252],ROW[251],ROW[250],ROW[249],ROW[248],ROW[247],ROW[246],ROW[245],ROW[244],ROW[243],ROW[242],ROW[241],ROW[240],ROW[239],ROW[238],ROW[237],ROW[236],ROW[235],ROW[234],ROW[233],ROW[232],ROW[231],ROW[230],ROW[229],ROW[228],ROW[227],ROW[226],ROW[225],ROW[224],ROW[223],ROW[222],ROW[221],ROW[220],ROW[219],ROW[218],ROW[217],ROW[216],ROW[215],ROW[214],ROW[213],ROW[212],ROW[211],ROW[210],ROW[209],ROW[208],ROW[207],ROW[206],ROW[205],ROW[204],ROW[203],ROW[202],ROW[201],ROW[200],ROW[199],ROW[198],ROW[197],ROW[196],ROW[195],ROW[194],ROW[193],ROW[192],ROW[191],ROW[190],ROW[189],ROW[188],ROW[187],ROW[186],ROW[185],ROW[184],ROW[183],ROW[182],ROW[181],ROW[180],ROW[179],ROW[178],ROW[177],ROW[176],ROW[175],ROW[174],ROW[173],ROW[172],ROW[171],ROW[170],ROW[169],ROW[168],ROW[167],ROW[166],ROW[165],ROW[164],ROW[163],ROW[162],ROW[161],ROW[160],ROW[159],ROW[158],ROW[157],ROW[156],ROW[155],ROW[154],ROW[153],ROW[152],ROW[151],ROW[150],ROW[149],ROW[148],ROW[147],ROW[146],ROW[145],ROW[144],ROW[143],ROW[142],ROW[141],ROW[140],ROW[139],ROW[138],ROW[137],ROW[136],ROW[135],ROW[134],ROW[133],ROW[132],ROW[131],ROW[130],ROW[129],ROW[128],ROW[127],ROW[126],ROW[125],ROW[124],ROW[123],ROW[122],ROW[121],ROW[120],ROW[119],ROW[118],ROW[117],ROW[116],ROW[115],ROW[114],ROW[113],ROW[112],ROW[111],ROW[110],ROW[109],ROW[108],ROW[107],ROW[106],ROW[105],ROW[104],ROW[103],ROW[102],ROW[101],ROW[100],ROW[99],ROW[98],ROW[97],ROW[96],ROW[95],ROW[94],ROW[93],ROW[92],ROW[91],ROW[90],ROW[89],ROW[88],ROW[87],ROW[86],ROW[85],ROW[84],ROW[83],ROW[82],ROW[81],ROW[80],ROW[79],ROW[78],ROW[77],ROW[76],ROW[75],ROW[74],ROW[73],ROW[72],ROW[71],ROW[70],ROW[69],ROW[68],ROW[67],ROW[66],ROW[65],ROW[64],ROW[63],ROW[62],ROW[61],ROW[60],ROW[59],ROW[58],ROW[57],ROW[56],ROW[55],ROW[54],ROW[53],ROW[52],ROW[51],ROW[50],ROW[49],ROW[48],ROW[47],ROW[46],ROW[45],ROW[44],ROW[43],ROW[42],ROW[41],ROW[40],ROW[39],ROW[38],ROW[37],ROW[36],ROW[35],ROW[34],ROW[33],ROW[32],ROW[31],ROW[30],ROW[29],ROW[28],ROW[27],ROW[26],ROW[25],ROW[24],ROW[23],ROW[22],ROW[21],ROW[20],ROW[19],ROW[18],ROW[17],ROW[16],ROW[15],ROW[14],ROW[13],ROW[12],ROW[11],ROW[10],ROW[9],ROW[8],ROW[7],ROW[6],ROW[5],ROW[4],ROW[3],ROW[2],ROW[1],ROW[0] COL[3],COL[2],COL[1],COL[0]
*.ipin A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2]
*.opin
*+ ROW[255],ROW[254],ROW[253],ROW[252],ROW[251],ROW[250],ROW[249],ROW[248],ROW[247],ROW[246],ROW[245],ROW[244],ROW[243],ROW[242],ROW[241],ROW[240],ROW[239],ROW[238],ROW[237],ROW[236],ROW[235],ROW[234],ROW[233],ROW[232],ROW[231],ROW[230],ROW[229],ROW[228],ROW[227],ROW[226],ROW[225],ROW[224],ROW[223],ROW[222],ROW[221],ROW[220],ROW[219],ROW[218],ROW[217],ROW[216],ROW[215],ROW[214],ROW[213],ROW[212],ROW[211],ROW[210],ROW[209],ROW[208],ROW[207],ROW[206],ROW[205],ROW[204],ROW[203],ROW[202],ROW[201],ROW[200],ROW[199],ROW[198],ROW[197],ROW[196],ROW[195],ROW[194],ROW[193],ROW[192],ROW[191],ROW[190],ROW[189],ROW[188],ROW[187],ROW[186],ROW[185],ROW[184],ROW[183],ROW[182],ROW[181],ROW[180],ROW[179],ROW[178],ROW[177],ROW[176],ROW[175],ROW[174],ROW[173],ROW[172],ROW[171],ROW[170],ROW[169],ROW[168],ROW[167],ROW[166],ROW[165],ROW[164],ROW[163],ROW[162],ROW[161],ROW[160],ROW[159],ROW[158],ROW[157],ROW[156],ROW[155],ROW[154],ROW[153],ROW[152],ROW[151],ROW[150],ROW[149],ROW[148],ROW[147],ROW[146],ROW[145],ROW[144],ROW[143],ROW[142],ROW[141],ROW[140],ROW[139],ROW[138],ROW[137],ROW[136],ROW[135],ROW[134],ROW[133],ROW[132],ROW[131],ROW[130],ROW[129],ROW[128],ROW[127],ROW[126],ROW[125],ROW[124],ROW[123],ROW[122],ROW[121],ROW[120],ROW[119],ROW[118],ROW[117],ROW[116],ROW[115],ROW[114],ROW[113],ROW[112],ROW[111],ROW[110],ROW[109],ROW[108],ROW[107],ROW[106],ROW[105],ROW[104],ROW[103],ROW[102],ROW[101],ROW[100],ROW[99],ROW[98],ROW[97],ROW[96],ROW[95],ROW[94],ROW[93],ROW[92],ROW[91],ROW[90],ROW[89],ROW[88],ROW[87],ROW[86],ROW[85],ROW[84],ROW[83],ROW[82],ROW[81],ROW[80],ROW[79],ROW[78],ROW[77],ROW[76],ROW[75],ROW[74],ROW[73],ROW[72],ROW[71],ROW[70],ROW[69],ROW[68],ROW[67],ROW[66],ROW[65],ROW[64],ROW[63],ROW[62],ROW[61],ROW[60],ROW[59],ROW[58],ROW[57],ROW[56],ROW[55],ROW[54],ROW[53],ROW[52],ROW[51],ROW[50],ROW[49],ROW[48],ROW[47],ROW[46],ROW[45],ROW[44],ROW[43],ROW[42],ROW[41],ROW[40],ROW[39],ROW[38],ROW[37],ROW[36],ROW[35],ROW[34],ROW[33],ROW[32],ROW[31],ROW[30],ROW[29],ROW[28],ROW[27],ROW[26],ROW[25],ROW[24],ROW[23],ROW[22],ROW[21],ROW[20],ROW[19],ROW[18],ROW[17],ROW[16],ROW[15],ROW[14],ROW[13],ROW[12],ROW[11],ROW[10],ROW[9],ROW[8],ROW[7],ROW[6],ROW[5],ROW[4],ROW[3],ROW[2],ROW[1],ROW[0]
*.opin COL[3],COL[2],COL[1],COL[0]
x1 A[11] A[10] A[9] A[8] SEL_hi[15] SEL_hi[14] SEL_hi[13] SEL_hi[12] SEL_hi[11] SEL_hi[10] SEL_hi[9]
+ SEL_hi[8] SEL_hi[7] SEL_hi[6] SEL_hi[5] SEL_hi[4] SEL_hi[3] SEL_hi[2] SEL_hi[1] SEL_hi[0] rom_dec_4b
x3 A[3] A[2] net9[3] net9[2] net9[1] net9[0] rom_dec_2b
x2 A[7] A[6] A[5] A[4] SEL_lo[15] SEL_lo[14] SEL_lo[13] SEL_lo[12] SEL_lo[11] SEL_lo[10] SEL_lo[9]
+ SEL_lo[8] SEL_lo[7] SEL_lo[6] SEL_lo[5] SEL_lo[4] SEL_lo[3] SEL_lo[2] SEL_lo[1] SEL_lo[0] rom_dec_4b
x1[3] net9[3] COL[3] not
x1[2] net9[2] COL[2] not
x1[1] net9[1] COL[1] not
x1[0] net9[0] COL[0] not
x5 net1[3] net1[2] net1[1] net1[0] ROW[31] ROW[30] ROW[29] ROW[28] ROW[27] ROW[26] ROW[25] ROW[24]
+ ROW[23] ROW[22] ROW[21] ROW[20] ROW[19] ROW[18] ROW[17] ROW[16] net2[3] net2[2] net2[1] net2[0]
+ rom_dec_cell
x6 net1[3] net1[2] net1[1] net1[0] ROW[47] ROW[46] ROW[45] ROW[44] ROW[43] ROW[42] ROW[41] ROW[40]
+ ROW[39] ROW[38] ROW[37] ROW[36] ROW[35] ROW[34] ROW[33] ROW[32] net3[3] net3[2] net3[1] net3[0]
+ rom_dec_cell
x7 net1[3] net1[2] net1[1] net1[0] ROW[15] ROW[14] ROW[13] ROW[12] ROW[11] ROW[10] ROW[9] ROW[8]
+ ROW[7] ROW[6] ROW[5] ROW[4] ROW[3] ROW[2] ROW[1] ROW[0] net4[3] net4[2] net4[1] net4[0] rom_dec_cell
x8 net1[3] net1[2] net1[1] net1[0] ROW[63] ROW[62] ROW[61] ROW[60] ROW[59] ROW[58] ROW[57] ROW[56]
+ ROW[55] ROW[54] ROW[53] ROW[52] ROW[51] ROW[50] ROW[49] ROW[48] net5[3] net5[2] net5[1] net5[0]
+ rom_dec_cell
x4 net6[3] net6[2] net6[1] net6[0] ROW[95] ROW[94] ROW[93] ROW[92] ROW[91] ROW[90] ROW[89] ROW[88]
+ ROW[87] ROW[86] ROW[85] ROW[84] ROW[83] ROW[82] ROW[81] ROW[80] net2[3] net2[2] net2[1] net2[0]
+ rom_dec_cell
x9 net6[3] net6[2] net6[1] net6[0] ROW[111] ROW[110] ROW[109] ROW[108] ROW[107] ROW[106] ROW[105]
+ ROW[104] ROW[103] ROW[102] ROW[101] ROW[100] ROW[99] ROW[98] ROW[97] ROW[96] net3[3] net3[2] net3[1] net3[0]
+ rom_dec_cell
x10 net6[3] net6[2] net6[1] net6[0] ROW[79] ROW[78] ROW[77] ROW[76] ROW[75] ROW[74] ROW[73] ROW[72]
+ ROW[71] ROW[70] ROW[69] ROW[68] ROW[67] ROW[66] ROW[65] ROW[64] net4[3] net4[2] net4[1] net4[0]
+ rom_dec_cell
x11 net6[3] net6[2] net6[1] net6[0] ROW[127] ROW[126] ROW[125] ROW[124] ROW[123] ROW[122] ROW[121]
+ ROW[120] ROW[119] ROW[118] ROW[117] ROW[116] ROW[115] ROW[114] ROW[113] ROW[112] net5[3] net5[2] net5[1]
+ net5[0] rom_dec_cell
x12 net7[3] net7[2] net7[1] net7[0] ROW[159] ROW[158] ROW[157] ROW[156] ROW[155] ROW[154] ROW[153]
+ ROW[152] ROW[151] ROW[150] ROW[149] ROW[148] ROW[147] ROW[146] ROW[145] ROW[144] net2[3] net2[2] net2[1]
+ net2[0] rom_dec_cell
x13 net7[3] net7[2] net7[1] net7[0] ROW[175] ROW[174] ROW[173] ROW[172] ROW[171] ROW[170] ROW[169]
+ ROW[168] ROW[167] ROW[166] ROW[165] ROW[164] ROW[163] ROW[162] ROW[161] ROW[160] net3[3] net3[2] net3[1]
+ net3[0] rom_dec_cell
x14 net7[3] net7[2] net7[1] net7[0] ROW[143] ROW[142] ROW[141] ROW[140] ROW[139] ROW[138] ROW[137]
+ ROW[136] ROW[135] ROW[134] ROW[133] ROW[132] ROW[131] ROW[130] ROW[129] ROW[128] net4[3] net4[2] net4[1]
+ net4[0] rom_dec_cell
x15 net7[3] net7[2] net7[1] net7[0] ROW[191] ROW[190] ROW[189] ROW[188] ROW[187] ROW[186] ROW[185]
+ ROW[184] ROW[183] ROW[182] ROW[181] ROW[180] ROW[179] ROW[178] ROW[177] ROW[176] net5[3] net5[2] net5[1]
+ net5[0] rom_dec_cell
x16 net8[3] net8[2] net8[1] net8[0] ROW[223] ROW[222] ROW[221] ROW[220] ROW[219] ROW[218] ROW[217]
+ ROW[216] ROW[215] ROW[214] ROW[213] ROW[212] ROW[211] ROW[210] ROW[209] ROW[208] net2[3] net2[2] net2[1]
+ net2[0] rom_dec_cell
x17 net8[3] net8[2] net8[1] net8[0] ROW[239] ROW[238] ROW[237] ROW[236] ROW[235] ROW[234] ROW[233]
+ ROW[232] ROW[231] ROW[230] ROW[229] ROW[228] ROW[227] ROW[226] ROW[225] ROW[224] net3[3] net3[2] net3[1]
+ net3[0] rom_dec_cell
x18 net8[3] net8[2] net8[1] net8[0] ROW[207] ROW[206] ROW[205] ROW[204] ROW[203] ROW[202] ROW[201]
+ ROW[200] ROW[199] ROW[198] ROW[197] ROW[196] ROW[195] ROW[194] ROW[193] ROW[192] net4[3] net4[2] net4[1]
+ net4[0] rom_dec_cell
x19 net8[3] net8[2] net8[1] net8[0] ROW[255] ROW[254] ROW[253] ROW[252] ROW[251] ROW[250] ROW[249]
+ ROW[248] ROW[247] ROW[246] ROW[245] ROW[244] ROW[243] ROW[242] ROW[241] ROW[240] net5[3] net5[2] net5[1]
+ net5[0] rom_dec_cell
x2[3] SEL_hi[15] net8[3] not
x2[2] SEL_hi[14] net8[2] not
x2[1] SEL_hi[13] net8[1] not
x2[0] SEL_hi[12] net8[0] not
x3[3] SEL_hi[11] net7[3] not
x3[2] SEL_hi[10] net7[2] not
x3[1] SEL_hi[9] net7[1] not
x3[0] SEL_hi[8] net7[0] not
x4[3] SEL_hi[7] net6[3] not
x4[2] SEL_hi[6] net6[2] not
x4[1] SEL_hi[5] net6[1] not
x4[0] SEL_hi[4] net6[0] not
x5[3] SEL_hi[3] net1[3] not
x5[2] SEL_hi[2] net1[2] not
x5[1] SEL_hi[1] net1[1] not
x5[0] SEL_hi[0] net1[0] not
x6[3] SEL_lo[3] net4[3] not
x6[2] SEL_lo[2] net4[2] not
x6[1] SEL_lo[1] net4[1] not
x6[0] SEL_lo[0] net4[0] not
x7[3] SEL_lo[7] net2[3] not
x7[2] SEL_lo[6] net2[2] not
x7[1] SEL_lo[5] net2[1] not
x7[0] SEL_lo[4] net2[0] not
x8[3] SEL_lo[11] net3[3] not
x8[2] SEL_lo[10] net3[2] not
x8[1] SEL_lo[9] net3[1] not
x8[0] SEL_lo[8] net3[0] not
x9[3] SEL_lo[15] net5[3] not
x9[2] SEL_lo[14] net5[2] not
x9[1] SEL_lo[13] net5[1] not
x9[0] SEL_lo[12] net5[0] not
**.ends

* expanding   symbol:  rom_dec_4b.sym # of pins=2
** sym_path: /media/FlexRV32/asic/blocks/rom/rom_dec_4b.sym
** sch_path: /media/FlexRV32/asic/blocks/rom/rom_dec_4b.sch
.subckt rom_dec_4b A[3] A[2] A[1] A[0] SEL[15] SEL[14] SEL[13] SEL[12] SEL[11] SEL[10] SEL[9] SEL[8]
+ SEL[7] SEL[6] SEL[5] SEL[4] SEL[3] SEL[2] SEL[1] SEL[0]
*.opin
*+ SEL[15],SEL[14],SEL[13],SEL[12],SEL[11],SEL[10],SEL[9],SEL[8],SEL[7],SEL[6],SEL[5],SEL[4],SEL[3],SEL[2],SEL[1],SEL[0]
*.ipin A[3],A[2],A[1],A[0]
x1 A[1] A[0] SEL_lo[3] SEL_lo[2] SEL_lo[1] SEL_lo[0] rom_dec_2b
x2 A[3] A[2] SEL_hi[3] SEL_hi[2] SEL_hi[1] SEL_hi[0] rom_dec_2b
x4 SEL_hi[0] SEL_lo[1] SEL[1] rom_nor2
x3 SEL_hi[0] SEL_lo[0] SEL[0] rom_nor2
x6 SEL_hi[0] SEL_lo[3] SEL[3] rom_nor2
x5 SEL_hi[0] SEL_lo[2] SEL[2] rom_nor2
x7 SEL_hi[1] SEL_lo[1] SEL[5] rom_nor2
x8 SEL_hi[1] SEL_lo[0] SEL[4] rom_nor2
x9 SEL_hi[1] SEL_lo[3] SEL[7] rom_nor2
x10 SEL_hi[1] SEL_lo[2] SEL[6] rom_nor2
x11 SEL_hi[2] SEL_lo[1] SEL[9] rom_nor2
x12 SEL_hi[2] SEL_lo[0] SEL[8] rom_nor2
x13 SEL_hi[2] SEL_lo[3] SEL[11] rom_nor2
x14 SEL_hi[2] SEL_lo[2] SEL[10] rom_nor2
x15 SEL_hi[3] SEL_lo[1] SEL[13] rom_nor2
x16 SEL_hi[3] SEL_lo[0] SEL[12] rom_nor2
x17 SEL_hi[3] SEL_lo[3] SEL[15] rom_nor2
x18 SEL_hi[3] SEL_lo[2] SEL[14] rom_nor2
.ends


* expanding   symbol:  rom_dec_2b.sym # of pins=2
** sym_path: /media/FlexRV32/asic/blocks/rom/rom_dec_2b.sym
** sch_path: /media/FlexRV32/asic/blocks/rom/rom_dec_2b.sch
.subckt rom_dec_2b A[1] A[0] SEL_n[3] SEL_n[2] SEL_n[1] SEL_n[0]
*.ipin A[1],A[0]
*.opin SEL_n[3],SEL_n[2],SEL_n[1],SEL_n[0]
x1 SEL_n[0] net1 net3 rom_nand2
x2 SEL_n[1] net2 net3 rom_nand2
x3 SEL_n[2] net1 net4 rom_nand2
x4 SEL_n[3] net2 net4 rom_nand2
x5 A[0] net1 not
x6 A[1] net3 not
x7 net1 net2 not
x8 net3 net4 not
.ends


* expanding   symbol:  ../../elements/logic/not.sym # of pins=2
** sym_path: /media/FlexRV32/asic/elements/logic/not.sym
** sch_path: /media/FlexRV32/asic/elements/logic/not.sch
.subckt not A Y
*.ipin A
*.opin Y
XM1 Y A VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
.ends


* expanding   symbol:  rom_dec_cell.sym # of pins=3
** sym_path: /media/FlexRV32/asic/blocks/rom/rom_dec_cell.sym
** sch_path: /media/FlexRV32/asic/blocks/rom/rom_dec_cell.sch
.subckt rom_dec_cell ROW[3] ROW[2] ROW[1] ROW[0] SEL[15] SEL[14] SEL[13] SEL[12] SEL[11] SEL[10]
+ SEL[9] SEL[8] SEL[7] SEL[6] SEL[5] SEL[4] SEL[3] SEL[2] SEL[1] SEL[0] COL[3] COL[2] COL[1] COL[0]
*.opin
*+ SEL[15],SEL[14],SEL[13],SEL[12],SEL[11],SEL[10],SEL[9],SEL[8],SEL[7],SEL[6],SEL[5],SEL[4],SEL[3],SEL[2],SEL[1],SEL[0]
*.ipin ROW[3],ROW[2],ROW[1],ROW[0]
*.ipin COL[3],COL[2],COL[1],COL[0]
x1 ROW[0] net1 not
x2 ROW[1] net2 not
x3 ROW[2] net3 not
x4 ROW[3] net4 not
x5 COL[0] net5 not
x6 COL[1] net6 not
x7 COL[2] net7 not
x8 COL[3] net8 not
x9 SEL[0] net1 net5 rom_nand2
x10 SEL[4] net2 net5 rom_nand2
x11 SEL[8] net3 net5 rom_nand2
x12 SEL[12] net4 net5 rom_nand2
x13 SEL[1] net1 net6 rom_nand2
x14 SEL[5] net2 net6 rom_nand2
x15 SEL[9] net3 net6 rom_nand2
x16 SEL[13] net4 net6 rom_nand2
x17 SEL[2] net1 net7 rom_nand2
x18 SEL[6] net2 net7 rom_nand2
x19 SEL[10] net3 net7 rom_nand2
x20 SEL[14] net4 net7 rom_nand2
x21 SEL[3] net1 net8 rom_nand2
x22 SEL[7] net2 net8 rom_nand2
x23 SEL[11] net3 net8 rom_nand2
x24 SEL[15] net4 net8 rom_nand2
.ends


* expanding   symbol:  rom_nor2.sym # of pins=3
** sym_path: /media/FlexRV32/asic/blocks/rom/rom_nor2.sym
** sch_path: /media/FlexRV32/asic/blocks/rom/rom_nor2.sch
.subckt rom_nor2 A B NOR
*.ipin A
*.opin NOR
*.ipin B
XM4 net1 A VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM5 NOR B net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM9 NOR B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM10 NOR A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
.ends


* expanding   symbol:  ./rom_nand2.sym # of pins=3
** sym_path: /media/FlexRV32/asic/blocks/rom/rom_nand2.sym
** sch_path: /media/FlexRV32/asic/blocks/rom/rom_nand2.sch
.subckt rom_nand2 NAND A B
*.ipin A
*.opin NAND
*.ipin B
XM2 NAND B VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM3 NAND A VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM6 NAND A p0 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM7 p0 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
.ends

.GLOBAL VCC
.GLOBAL VSS
.end
